library ieee;
use ieee.std_logic_1164.all;

entity decoderInstru is
  port ( opcode : in std_logic_vector(5 downto 0);
         saida : out std_logic_vector(14 downto 0)
  );
end entity;

architecture comportamento of decoderInstru is

  constant LW  : std_logic_vector(5 downto 0) := "100011";
  constant SW  : std_logic_vector(5 downto 0) := "101011";
  constant BEQ : std_logic_vector(5 downto 0) := "000100";
  constant JMP : std_logic_vector(5 downto 0) := "000010";
  constant INST_R : std_logic_vector(5 downto 0) := "000000";
  

  begin

 
saida <=   "0011" & LW & "01010" when opcode = LW else
			  "0001" & SW & "00001" when opcode = SW else
			  "0000" & BEQ & "00100" when opcode = BEQ else
			  "1000" & JMP & "00000" when opcode = JMP else
			  "0110" & INST_R & "10000" when opcode = INST_R else
			  "000000000000000"; -- NOP para intrucoes indefinidas
end architecture;
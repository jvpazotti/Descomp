library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 13;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is
  
  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI	 : std_logic_vector(3 downto 0) := "0100";
  constant STA	 : std_logic_vector(3 downto 0) := "0101";
  constant JMP : std_logic_vector(3 downto 0) := "0110";
  constant JEQ : std_logic_vector(3 downto 0) := "0111";
  constant CEQ : std_logic_vector(3 downto 0) := "1000";
  constant JSR : std_logic_vector(3 downto 0) := "1001";
  constant RET : std_logic_vector(3 downto 0) := "1010";
  constant GT : std_logic_vector(3 downto 0) := "1011";
  constant JGT : std_logic_vector(3 downto 0) := "1100";
  
  constant R0:    std_logic_vector (1 DOWNTO 0)	:= "00";
  constant R1:    std_logic_vector (1 DOWNTO 0)	:= "01";
  constant R2:    std_logic_vector (1 DOWNTO 0)	:= "10";
  constant R3:    std_logic_vector (1 DOWNTO 0)	:= "11";


  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Reset_A, Operacao_ULA
      -- Inicializa os endereços:
tmp(0) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(1) := R0 & LDI  & '0' & x"00";	-- LDI R0, $0	#Início do Setup
tmp(2) := R0 & STA  & '1' & x"20";	-- STA R0, @288	#Zerando hexas
tmp(3) := R0 & STA  & '1' & x"21";	-- STA R0, @289
tmp(4) := R0 & STA  & '1' & x"22";	-- STA R0, @290
tmp(5) := R0 & STA  & '1' & x"23";	-- STA R0, @291
tmp(6) := R0 & STA  & '1' & x"24";	-- STA R0, @292
tmp(7) := R0 & STA  & '1' & x"25";	-- STA R0, @293
tmp(8) := R0 & STA  & '1' & x"00";	-- STA R0, @256	#Zerando leds
tmp(9) := R0 & STA  & '1' & x"01";	-- STA R0, @257
tmp(10) := R0 & STA  & '1' & x"02";	-- STA R0, @258
tmp(11) := R0 & STA  & '0' & x"00";	-- STA R0, @0	#Armazenando 0 em unidade, dezena, centena, etc
tmp(12) := R0 & STA  & '0' & x"01";	-- STA R0, @1
tmp(13) := R0 & STA  & '0' & x"02";	-- STA R0, @2
tmp(14) := R0 & STA  & '0' & x"03";	-- STA R0, @3
tmp(15) := R0 & STA  & '0' & x"04";	-- STA R0, @4
tmp(16) := R0 & STA  & '0' & x"05";	-- STA R0, @5
tmp(17) := R0 & STA  & '0' & x"06";	-- STA R0, @6	#Constante de comparacao (0)
tmp(18) := R0 & STA  & '0' & x"0F";	-- STA R0, @15	#Flag que para contagem
tmp(19) := R0 & STA  & '1' & x"FE";	-- STA R0, @510
tmp(20) := R0 & STA  & '1' & x"FF";	-- STA R0, @511
tmp(21) := R0 & STA  & '1' & x"FD";	-- STA R0, @509
tmp(22) := R0 & LDI  & '0' & x"01";	-- LDI R0, $1
tmp(23) := R0 & STA  & '0' & x"07";	-- STA R0, @7	#Constante de Incremento (1)
tmp(24) := R0 & LDI  & '0' & x"0A";	-- LDI R0, $10
tmp(25) := R0 & STA  & '0' & x"08";	-- STA R0, @8	#Constante de limite no display (10)
tmp(26) := R0 & LDI  & '0' & x"00";	-- LDI R0, $0
tmp(27) := R0 & STA  & '0' & x"09";	-- STA R0, @9	#Limite de contagem em unidade, dezena, centena, etc
tmp(28) := R0 & STA  & '0' & x"0A";	-- STA R0, @10
tmp(29) := R0 & STA  & '0' & x"0B";	-- STA R0, @11
tmp(30) := R0 & STA  & '0' & x"0C";	-- STA R0, @12
tmp(31) := R0 & STA  & '0' & x"0D";	-- STA R0, @13
tmp(32) := R0 & STA  & '0' & x"0E";	-- STA R0, @14
tmp(33) := R0 & LDI  & '0' & x"09";	-- LDI R0, $9
tmp(34) := R0 & STA  & '0' & x"10";	-- STA R0, @16	#Constante de limite de valor
tmp(35) := R0 & LDI  & '0' & x"05";	-- LDI R0, $5
tmp(36) := R0 & STA  & '0' & x"11";	-- STA R0, @17	#Constante de limite de valor de minutos e segundos
tmp(37) := R0 & LDI  & '0' & x"03";	-- LDI R0, $3
tmp(38) := R0 & STA  & '0' & x"12";	-- STA R0, @18	#Constante de limite de valor de horas1
tmp(39) := R0 & LDI  & '0' & x"02";	-- LDI R0, $2
tmp(40) := R0 & STA  & '0' & x"13";	-- STA R0, @19	#Constante de limite de valor de horas2
tmp(41) := R0 & LDI  & '0' & x"06";	-- LDI R0, $6
tmp(42) := R0 & STA  & '0' & x"14";	-- STA R0, @20
tmp(43) := R0 & LDI  & '0' & x"04";	-- LDI R0, $4
tmp(44) := R0 & STA  & '0' & x"15";	-- STA R0, @21
tmp(45) := R0 & NOP  & '0' & x"00";	-- NOP	#Loop principal
tmp(46) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	# Le o valor de KEY1
tmp(47) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	# Compara o valor de KEY1 com 0
tmp(48) := R0 & JEQ  & '0' & x"2D";	-- JEQ @INICIOLOOP	# Se for igual a 0, fica no aguardo para quando for 1
tmp(49) := R0 & JSR  & '0' & x"48";	-- JSR @CONFIGLIMITE	# Se for diferente de 0, entra na sub rotina de configuracao de Limite
tmp(50) := R0 & LDA  & '0' & x"06";	-- LDA R0, @6	#Carrega 0 no acumulador
tmp(51) := R0 & STA  & '1' & x"20";	-- STA R0, @288	# Zera o HEX1
tmp(52) := R0 & STA  & '1' & x"21";	-- STA R0, @289	# Zera o HEX2
tmp(53) := R0 & STA  & '1' & x"22";	-- STA R0, @290	# Zera o HEX3
tmp(54) := R0 & STA  & '1' & x"23";	-- STA R0, @291	# Zera o HEX4
tmp(55) := R0 & STA  & '1' & x"24";	-- STA R0, @292	# Zera o HEX5
tmp(56) := R0 & STA  & '1' & x"25";	-- STA R0, @293	# Zera o HEX6
tmp(57) := R0 & STA  & '1' & x"00";	-- STA R0, @256	# Zera os LEDS(7~0)
tmp(58) := R0 & STA  & '1' & x"02";	-- STA R0, @258	# Zera os LED(9)
tmp(59) := R0 & STA  & '1' & x"01";	-- STA R0, @257	# Zera os LED(8) 
tmp(60) := R0 & NOP  & '0' & x"00";	-- NOP	# Incrementa ate chegar no limite de contagem
tmp(61) := R2 & LDA  & '1' & x"60";	-- LDA R2, @352	# Le o valor de KEY0
tmp(62) := R2 & CEQ  & '0' & x"06";	-- CEQ R2, @6	# Compara o valor de KEY0 com 0
tmp(63) := R0 & JEQ  & '0' & x"41";	-- JEQ @PULA1	# Se for igual a 0, nao incrementa e atualiza os displays
tmp(64) := R0 & JSR  & '0' & x"F3";	-- JSR @INCREMENTA	# Se for diferente de 0, entra na sub rotina de incremento
tmp(65) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(66) := R0 & JSR  & '1' & x"30";	-- JSR @ATUALIZA	# Atualiza os displays
tmp(67) := R0 & JSR  & '1' & x"3E";	-- JSR @CHECALIMITE	# Checa pra ver se passou do limite setado
tmp(68) := R2 & LDA  & '0' & x"0F";	-- LDA R2, @15	# Le o valor da flag de inibir contagem
tmp(69) := R2 & CEQ  & '0' & x"06";	-- CEQ R2, @6	# Compara com 0 a flag (flag com valor 1 -> ativa, flag com valor 0 -> desativada)
tmp(70) := R0 & JEQ  & '0' & x"3C";	-- JEQ @INCREMENTADOR	#Se a flag for 0, pode continuar incrementando
tmp(71) := R0 & JMP  & '1' & x"61";	-- JMP @TRAVA	# Se for 1, trava a contagem
tmp(72) := R0 & NOP  & '0' & x"00";	-- NOP	#Rotina de configuracao de limite
tmp(73) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1	# Carrega o valor 1
tmp(74) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota no endereco dos LEDS(7-0)
tmp(75) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Limpa a leitura de KEY1
tmp(76) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(77) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(78) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(79) := R0 & JGT  & '0' & x"51";	-- JGT @VALORATUALIZADO	#Se for maior que 9, atualiza os displays
tmp(80) := R0 & JMP  & '0' & x"53";	-- JMP @IGNORA
tmp(81) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(82) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(83) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(84) := R1 & STA  & '1' & x"20";	-- STA R1, @288	# Hex 0
tmp(85) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	# Le KEY1
tmp(86) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara KEY1 com 0
tmp(87) := R0 & JEQ  & '0' & x"4C";	-- JEQ @ESPERAUNIDADE	#Se for 0, ou seja, nao esta apertado, espera ate apertar
tmp(88) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Limpa a leitura de KEY1
tmp(89) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(90) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(91) := R0 & JGT  & '0' & x"5D";	-- JGT @VALORATUALIZADO2	#Se for maior que 9, atualiza os displays
tmp(92) := R0 & JMP  & '0' & x"5F";	-- JMP @IGNORA2
tmp(93) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(94) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(95) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(96) := R1 & STA  & '0' & x"09";	-- STA R1, @9	#Armazena o valor das chaves no limite das unidades
tmp(97) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(98) := R1 & LDI  & '0' & x"04";	-- LDI R1, $4	#Carrega o valor 4
tmp(99) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(100) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(101) := R1 & GT  & '0' & x"11";	-- GT R1, @17	#Compara com 5
tmp(102) := R0 & JGT  & '0' & x"68";	-- JGT @VALORATUALIZADO3	#Se for maior que 5, atualiza os displays
tmp(103) := R0 & JMP  & '0' & x"6A";	-- JMP @IGNORA3
tmp(104) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(105) := R1 & LDI  & '0' & x"05";	-- LDI R1, $5
tmp(106) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(107) := R1 & STA  & '1' & x"21";	-- STA R1, @289	# Hex 1
tmp(108) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(109) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(110) := R0 & JEQ  & '0' & x"61";	-- JEQ @ESPERADEZENA	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(111) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(112) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(113) := R1 & GT  & '0' & x"11";	-- GT R1, @17	#Compara com 5
tmp(114) := R0 & JGT  & '0' & x"74";	-- JGT @VALORATUALIZADO4	#Se for maior que 5, atualiza os displays
tmp(115) := R0 & JMP  & '0' & x"76";	-- JMP @IGNORA4
tmp(116) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(117) := R1 & LDI  & '0' & x"05";	-- LDI R1, $5
tmp(118) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(119) := R1 & STA  & '0' & x"0A";	-- STA R1, @10	#Armazena o valor das chaves no limte das dezenas
tmp(120) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(121) := R1 & LDI  & '0' & x"10";	-- LDI R1, $16	# Carrega o valor 16 no acumulador
tmp(122) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(123) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(124) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(125) := R0 & JGT  & '0' & x"7F";	-- JGT @VALORATUALIZADO5	#Se for maior que 9, atualiza os displays
tmp(126) := R0 & JMP  & '0' & x"81";	-- JMP @IGNORA5
tmp(127) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(128) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(129) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(130) := R1 & STA  & '1' & x"22";	-- STA R1, @290	# Hex 2
tmp(131) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(132) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(133) := R0 & JEQ  & '0' & x"78";	-- JEQ @ESPERACENTENA	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(134) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(135) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(136) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(137) := R0 & JGT  & '0' & x"8B";	-- JGT @VALORATUALIZADO6	#Se for maior que 9, atualiza os displays
tmp(138) := R0 & JMP  & '0' & x"8D";	-- JMP @IGNORA6
tmp(139) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(140) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(141) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(142) := R1 & STA  & '0' & x"0B";	-- STA R1, @11	#Armazena o valor das chaves no limite das centenas
tmp(143) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(144) := R1 & LDI  & '0' & x"20";	-- LDI R1, $32	# Carrega o valor 32 no acumulador
tmp(145) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(146) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(147) := R1 & GT  & '0' & x"11";	-- GT R1, @17	#Compara com 5
tmp(148) := R0 & JGT  & '0' & x"96";	-- JGT @VALORATUALIZADO7	#Se for maior que 5, atualiza os displays
tmp(149) := R0 & JMP  & '0' & x"98";	-- JMP @IGNORA7
tmp(150) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(151) := R1 & LDI  & '0' & x"05";	-- LDI R1, $5
tmp(152) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(153) := R1 & STA  & '1' & x"23";	-- STA R1, @291	# Hex 3
tmp(154) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(155) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1
tmp(156) := R0 & JEQ  & '0' & x"8F";	-- JEQ @ESPERAUNIDADEMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(157) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(158) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(159) := R1 & GT  & '0' & x"11";	-- GT R1, @17	#Compara com 5
tmp(160) := R0 & JGT  & '0' & x"A2";	-- JGT @VALORATUALIZADO8	#Se for maior que 5, atualiza os displays
tmp(161) := R0 & JMP  & '0' & x"A4";	-- JMP @IGNORA8
tmp(162) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(163) := R1 & LDI  & '0' & x"05";	-- LDI R1, $5
tmp(164) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(165) := R1 & STA  & '0' & x"0C";	-- STA R1, @12	#Armazena o valor das chaves no limite das unidades de milhar
tmp(166) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(167) := R1 & LDI  & '0' & x"80";	-- LDI R1, $128	# Carrega o valor 128 no acumulador
tmp(168) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(169) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(170) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(171) := R0 & JGT  & '0' & x"AD";	-- JGT @VALORATUALIZADO9	#Se for maior que 9, atualiza os displays
tmp(172) := R0 & JMP  & '0' & x"AF";	-- JMP @IGNORA9
tmp(173) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(174) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(175) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(176) := R1 & STA  & '1' & x"24";	-- STA R1, @292	# Hex 4
tmp(177) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(178) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(179) := R0 & JEQ  & '0' & x"A6";	-- JEQ @ESPERADEZENAMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(180) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(181) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(182) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(183) := R0 & JGT  & '0' & x"B9";	-- JGT @VALORATUALIZADO10	#Se for maior que 9, atualiza os displays
tmp(184) := R0 & JMP  & '0' & x"BB";	-- JMP @IGNORA10
tmp(185) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(186) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(187) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(188) := R1 & STA  & '0' & x"0D";	-- STA R1, @13	#Armazena o valor das chaves no limite das dezenas de milhar
tmp(189) := R0 & JMP  & '0' & x"D5";	-- JMP @ESPERACENTENAMILHAR
tmp(190) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(191) := R1 & LDI  & '0' & x"80";	-- LDI R1, $128	# Carrega o valor 128 no acumulador
tmp(192) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(193) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(194) := R1 & GT  & '0' & x"12";	-- GT R1, @18	#Compara com 3
tmp(195) := R0 & JGT  & '0' & x"C5";	-- JGT @VALORATUALIZADO13	#Se for maior que 3, atualiza os displays
tmp(196) := R0 & JMP  & '0' & x"C7";	-- JMP @IGNORA13
tmp(197) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(198) := R1 & LDI  & '0' & x"03";	-- LDI R1, $3
tmp(199) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(200) := R1 & STA  & '1' & x"24";	-- STA R1, @292	# Hex 4
tmp(201) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(202) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(203) := R0 & JEQ  & '0' & x"BE";	-- JEQ @VOLTADEZENAMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(204) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(205) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(206) := R1 & GT  & '0' & x"12";	-- GT R1, @18	#Compara com 3
tmp(207) := R0 & JGT  & '0' & x"D1";	-- JGT @VALORATUALIZADO14	#Se for maior que 3, atualiza os displays
tmp(208) := R0 & JMP  & '0' & x"D3";	-- JMP @IGNORA14
tmp(209) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(210) := R1 & LDI  & '0' & x"03";	-- LDI R1, $3
tmp(211) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(212) := R1 & STA  & '0' & x"0D";	-- STA R1, @13	#Armazena o valor das chaves no limite das dezenas de milhar
tmp(213) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(214) := R1 & LDA  & '0' & x"06";	-- LDA R1, @6	#Carrega 0 no acumulador
tmp(215) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Zera o valor nos LEDS(7~0)
tmp(216) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1	# Carrega o valor 1 no acumulador
tmp(217) := R1 & STA  & '1' & x"01";	-- STA R1, @257	# Bota o valor nos LEDS
tmp(218) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(219) := R1 & GT  & '0' & x"13";	-- GT R1, @19	#Compara com 2
tmp(220) := R0 & JGT  & '0' & x"DE";	-- JGT @VALORATUALIZADO11	#Se for maior que 2, atualiza os displays
tmp(221) := R0 & JMP  & '0' & x"E0";	-- JMP @IGNORA11
tmp(222) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(223) := R1 & LDI  & '0' & x"02";	-- LDI R1, $2
tmp(224) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(225) := R1 & STA  & '1' & x"25";	-- STA R1, @293	# Hex 5
tmp(226) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(227) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1
tmp(228) := R0 & JEQ  & '0' & x"D5";	-- JEQ @ESPERACENTENAMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(229) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(230) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(231) := R1 & GT  & '0' & x"13";	-- GT R1, @19	#Compara com 2
tmp(232) := R0 & JGT  & '0' & x"EA";	-- JGT @VALORATUALIZADO12	#Se for maior que 2, atualiza os displays
tmp(233) := R0 & JMP  & '0' & x"EC";	-- JMP @IGNORA12
tmp(234) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(235) := R1 & LDI  & '0' & x"02";	-- LDI R1, $2
tmp(236) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(237) := R1 & STA  & '0' & x"0E";	-- STA R1, @14	#Armazena o valor das chaves no limite das centenas de milhar
tmp(238) := R1 & LDA  & '0' & x"0E";	-- LDA R1, @14
tmp(239) := R1 & SOMA  & '0' & x"0D";	-- SOMA R1, @13
tmp(240) := R1 & GT  & '0' & x"14";	-- GT R1, @20
tmp(241) := R0 & JGT  & '0' & x"BE";	-- JGT @VOLTADEZENAMILHAR
tmp(242) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(243) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(244) := R2 & STA  & '1' & x"FF";	-- STA R2, @511	#Limpa a leitura de KEY1
tmp(245) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(246) := R2 & LDA  & '0' & x"00";	-- LDA R2, @0	#Carrega o valor da unidade no acumulador
tmp(247) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na unidade
tmp(248) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara unidade com 10
tmp(249) := R0 & JEQ  & '0' & x"FC";	-- JEQ @UNIDADEPASSOU	#Se for igual a 10, incrementa a dezena
tmp(250) := R2 & STA  & '0' & x"00";	-- STA R2, @0	#Se for diferente de 10, armazena o valor da unidade
tmp(251) := R0 & RET  & '0' & x"00";	-- RET 	#Retorna para o LOOP principal
tmp(252) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(253) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(254) := R2 & STA  & '0' & x"00";	-- STA R2, @0	#Zera a unidade
tmp(255) := R2 & LDA  & '0' & x"01";	-- LDA R2, @1	#Carrega o valor da dezena no acumulador
tmp(256) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na dezena 
tmp(257) := R2 & CEQ  & '0' & x"11";	-- CEQ R2, @17	#Compara dezena com 6
tmp(258) := R2 & JEQ  & '1' & x"05";	-- JEQ R2, @DEZENAPASSOU	#Se for igual a 6, incrementa a centena
tmp(259) := R2 & STA  & '0' & x"01";	-- STA R2, @1	#Se for diferente de 6, armazena o valor da dezena
tmp(260) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(261) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(262) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(263) := R2 & STA  & '0' & x"01";	-- STA R2, @1	#Zera a dezena
tmp(264) := R2 & LDA  & '0' & x"02";	-- LDA R2, @2	#Carrega o valor da centena no acumulador
tmp(265) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na centena
tmp(266) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara centena com 10
tmp(267) := R0 & JEQ  & '1' & x"0E";	-- JEQ @CENTENAPASSOU	#Se for igual a 10, incrementa a unidade de milhar
tmp(268) := R2 & STA  & '0' & x"02";	-- STA R2, @2	#Se for diferente de 10, armazena o valor da centena
tmp(269) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(270) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(271) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(272) := R2 & STA  & '0' & x"02";	-- STA R2, @2	#Zera a centena
tmp(273) := R2 & LDA  & '0' & x"03";	-- LDA R2, @3	#Carrega o valor da unidade de milhar no acumulador
tmp(274) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na unidade de milhar
tmp(275) := R2 & CEQ  & '0' & x"11";	-- CEQ R2, @17	#Compara unidade de milhar com 6
tmp(276) := R0 & JEQ  & '1' & x"17";	-- JEQ @UNIDADEMILHARPASSOU	#Se for igual a 6, incrementa a dezena de milhar
tmp(277) := R2 & STA  & '0' & x"03";	-- STA R2, @3	#Se for diferente de 6, armazena o valor da unidade de milhar
tmp(278) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(279) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(280) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(281) := R2 & STA  & '0' & x"03";	-- STA R2, @3	#Zera a unidade de milhar
tmp(282) := R2 & LDA  & '0' & x"04";	-- LDA R2, @4	#Carrega o valor da dezena de milhar no acumulador
tmp(283) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na dezena de milhar
tmp(284) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara dezena de milhar com 10
tmp(285) := R0 & JEQ  & '1' & x"20";	-- JEQ @DEZENAMILHARPASSOU	#Se for igual a 10, incrementa a centena de milhar
tmp(286) := R2 & STA  & '0' & x"04";	-- STA R2, @4	#Se for diferente de 10, armazena o valor da dezena de milhar
tmp(287) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(288) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(289) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(290) := R2 & STA  & '0' & x"04";	-- STA R2, @4	#Zera a dezena de milhar
tmp(291) := R2 & LDA  & '0' & x"05";	-- LDA R2, @5	#Carrega o valor da centena de milhar no acumulador
tmp(292) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na centena de milhar
tmp(293) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara centena de milhar com 10
tmp(294) := R0 & JEQ  & '1' & x"29";	-- JEQ @CENTENAMILHARPASSOU	#Se for igual a 10, incrementa a unidade de milhao
tmp(295) := R2 & STA  & '0' & x"05";	-- STA R2, @5	#Se for diferente de 10, armazena o valor da centena de milhar
tmp(296) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(297) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(298) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(299) := R2 & STA  & '0' & x"05";	-- STA R2, @5	#Zera a centena de milhar
tmp(300) := R2 & LDI  & '0' & x"01";	-- LDI R2, $1	#Carrega 1 no acumulador
tmp(301) := R2 & STA  & '1' & x"02";	-- STA R2, @258	#Acende o LED(9)
tmp(302) := R2 & STA  & '0' & x"0F";	-- STA R2, @15	#Ativa a flag de inibir incremento
tmp(303) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(304) := R0 & NOP  & '0' & x"00";	-- NOP	#Atualiza os valores dos HEX
tmp(305) := R3 & LDA  & '0' & x"00";	-- LDA R3, @0	#Le o valor das unidades
tmp(306) := R3 & STA  & '1' & x"20";	-- STA R3, @288	#Armazena o valor das unidades no HEX0
tmp(307) := R3 & LDA  & '0' & x"01";	-- LDA R3, @1	#Le o valor das dezenas
tmp(308) := R3 & STA  & '1' & x"21";	-- STA R3, @289	#Armazena o valor das dezenas no HEX1
tmp(309) := R3 & LDA  & '0' & x"02";	-- LDA R3, @2	#Le o valor das centenas
tmp(310) := R3 & STA  & '1' & x"22";	-- STA R3, @290	#Armazena o valor das centenas no HEX2
tmp(311) := R3 & LDA  & '0' & x"03";	-- LDA R3, @3	#Le o valor das unidades de milhar
tmp(312) := R3 & STA  & '1' & x"23";	-- STA R3, @291	#Armazena o valor das unidades de milhar no HEX3
tmp(313) := R3 & LDA  & '0' & x"04";	-- LDA R3, @4	#Le o valor das dezenas de milhar
tmp(314) := R3 & STA  & '1' & x"24";	-- STA R3, @292	#Armazena o valor das dezenas de milhar no HEX4
tmp(315) := R3 & LDA  & '0' & x"05";	-- LDA R3, @5	#Le o valor das centenas de milhar
tmp(316) := R3 & STA  & '1' & x"25";	-- STA R3, @293	#Armazena o valor das centenas de milhar no HEX5
tmp(317) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(318) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(319) := R1 & LDA  & '0' & x"00";	-- LDA R1, @0	#Le o valor das unidades
tmp(320) := R1 & CEQ  & '0' & x"09";	-- CEQ R1, @9	#Compara com o valor limite das unidades
tmp(321) := R0 & JEQ  & '1' & x"43";	-- JEQ @CHECADEZENA	#Se for igual, checa se ocorre com as dezenas
tmp(322) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(323) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(324) := R1 & LDA  & '0' & x"01";	-- LDA R1, @1	#Le o valor das dezenas
tmp(325) := R1 & CEQ  & '0' & x"0A";	-- CEQ R1, @10	#Compara com o valor limite das dezenas
tmp(326) := R0 & JEQ  & '1' & x"48";	-- JEQ @CHECACENTENA	#Se for igual, checa se ocorre com as centenas
tmp(327) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(328) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(329) := R1 & LDA  & '0' & x"02";	-- LDA R1, @2	#Le o valor das centenas
tmp(330) := R1 & CEQ  & '0' & x"0B";	-- CEQ R1, @11	#Compara com o valor limite das centenas
tmp(331) := R0 & JEQ  & '1' & x"4D";	-- JEQ @CHECAUNIDADEMILHAR	#Se for igual, checa se ocorre com as unidades de milhar
tmp(332) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(333) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(334) := R1 & LDA  & '0' & x"03";	-- LDA R1, @3	# Le o valor das unidades de milhar
tmp(335) := R1 & CEQ  & '0' & x"0C";	-- CEQ R1, @12	# Compara com o valor limite das unidades de milhar 
tmp(336) := R0 & JEQ  & '1' & x"52";	-- JEQ @CHECADEZENAMILHAR	#Se for igual, checa se ocorre com as dezenas de milhar
tmp(337) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(338) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(339) := R1 & LDA  & '0' & x"04";	-- LDA R1, @4	# Le o valor das dezenas de milhar
tmp(340) := R1 & CEQ  & '0' & x"0D";	-- CEQ R1, @13	# Compara com o valor limite das dezenas de milhar 
tmp(341) := R0 & JEQ  & '1' & x"57";	-- JEQ @CHECACENTENAMILHAR	#Se for igual, checa se ocorre com as centenas de milhar
tmp(342) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(343) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(344) := R1 & LDA  & '0' & x"05";	-- LDA R1, @5	# Le o valor das centenas de milhar
tmp(345) := R1 & CEQ  & '0' & x"0E";	-- CEQ R1, @14	# Compara com o valor limite das centenas de milhar 
tmp(346) := R0 & JEQ  & '1' & x"5C";	-- JEQ @BATEUNOLIMITE	#Se for igual, indica que o limite foi batido
tmp(347) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(348) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(349) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1	#Atribui o valor 1 no acumulador
tmp(350) := R1 & STA  & '0' & x"0F";	-- STA R1, @15	#Ativa a flag de parar contagem
tmp(351) := R1 & STA  & '1' & x"02";	-- STA R1, @258	#Ativa o LED de limite atingido 
tmp(352) := R0 & RET  & '0' & x"00";	-- RET	#Retorna pro LOOP principal
tmp(353) := R0 & NOP  & '0' & x"00";	-- NOP	#Trava a contagem
tmp(354) := R3 & LDI  & '0' & x"01";	-- LDI R3, $1
tmp(355) := R3 & STA  & '1' & x"00";	-- STA R3, @256
tmp(356) := R3 & LDA  & '1' & x"64";	-- LDA R3, @356	#Le o valor do botao FPGA
tmp(357) := R3 & CEQ  & '0' & x"06";	-- CEQ R3, @6	#Compara com 0 o botao FPGA
tmp(358) := R0 & JEQ  & '1' & x"61";	-- JEQ @TRAVA	#Se for igual, continua travado
tmp(359) := R0 & JMP  & '0' & x"00";	-- JMP @RESTART	#Se for diferente, reinicia a contagem




        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;
library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 13;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is
  
  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI	 : std_logic_vector(3 downto 0) := "0100";
  constant STA	 : std_logic_vector(3 downto 0) := "0101";
  constant JMP : std_logic_vector(3 downto 0) := "0110";
  constant JEQ : std_logic_vector(3 downto 0) := "0111";
  constant CEQ : std_logic_vector(3 downto 0) := "1000";
  constant JSR : std_logic_vector(3 downto 0) := "1001";
  constant RET : std_logic_vector(3 downto 0) := "1010";
  constant GT : std_logic_vector(3 downto 0) := "1011";
  constant JGT : std_logic_vector(3 downto 0) := "1100";
  
  constant R0:    std_logic_vector (1 DOWNTO 0)	:= "00";
  constant R1:    std_logic_vector (1 DOWNTO 0)	:= "01";
  constant R2:    std_logic_vector (1 DOWNTO 0)	:= "10";
  constant R3:    std_logic_vector (1 DOWNTO 0)	:= "11";


  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Reset_A, Operacao_ULA
      -- Inicializa os endereços:
tmp(0) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(1) := R0 & LDI  & '0' & x"00";	-- LDI R0, $0	#Início do Setup
tmp(2) := R0 & STA  & '1' & x"20";	-- STA R0, @288	#Zerando hexas
tmp(3) := R0 & STA  & '1' & x"21";	-- STA R0, @289
tmp(4) := R0 & STA  & '1' & x"22";	-- STA R0, @290
tmp(5) := R0 & STA  & '1' & x"23";	-- STA R0, @291
tmp(6) := R0 & STA  & '1' & x"24";	-- STA R0, @292
tmp(7) := R0 & STA  & '1' & x"25";	-- STA R0, @293
tmp(8) := R0 & STA  & '1' & x"00";	-- STA R0, @256	#Zerando leds
tmp(9) := R0 & STA  & '1' & x"01";	-- STA R0, @257
tmp(10) := R0 & STA  & '1' & x"02";	-- STA R0, @258
tmp(11) := R0 & STA  & '0' & x"00";	-- STA R0, @0	#Armazenando 0 em unidade, dezena, centena, etc
tmp(12) := R0 & STA  & '0' & x"01";	-- STA R0, @1
tmp(13) := R0 & STA  & '0' & x"02";	-- STA R0, @2
tmp(14) := R0 & STA  & '0' & x"03";	-- STA R0, @3
tmp(15) := R0 & STA  & '0' & x"04";	-- STA R0, @4
tmp(16) := R0 & STA  & '0' & x"05";	-- STA R0, @5
tmp(17) := R0 & STA  & '0' & x"06";	-- STA R0, @6	#Constante de comparacao (0)
tmp(18) := R0 & STA  & '1' & x"FE";	-- STA R0, @510
tmp(19) := R0 & STA  & '1' & x"FF";	-- STA R0, @511
tmp(20) := R0 & STA  & '1' & x"FD";	-- STA R0, @509
tmp(21) := R0 & LDI  & '0' & x"01";	-- LDI R0, $1
tmp(22) := R0 & STA  & '0' & x"07";	-- STA R0, @7	#Constante de Incremento (1)
tmp(23) := R0 & LDI  & '0' & x"0A";	-- LDI R0, $10
tmp(24) := R0 & STA  & '0' & x"08";	-- STA R0, @8	#Constante de limite no display (10)
tmp(25) := R0 & LDI  & '0' & x"00";	-- LDI R0, $0
tmp(26) := R0 & STA  & '0' & x"09";	-- STA R0, @9	#Limite de contagem em unidade, dezena, centena, etc
tmp(27) := R0 & STA  & '0' & x"0A";	-- STA R0, @10
tmp(28) := R0 & STA  & '0' & x"0B";	-- STA R0, @11
tmp(29) := R0 & STA  & '0' & x"0C";	-- STA R0, @12
tmp(30) := R0 & STA  & '0' & x"0D";	-- STA R0, @13
tmp(31) := R0 & STA  & '0' & x"0E";	-- STA R0, @14
tmp(32) := R0 & STA  & '0' & x"0F";	-- STA R0, @15
tmp(33) := R0 & LDI  & '0' & x"09";	-- LDI R0, $9
tmp(34) := R0 & STA  & '0' & x"10";	-- STA R0, @16	#Constante de limite de valor(9)
tmp(35) := R0 & LDI  & '0' & x"05";	-- LDI R0, $5
tmp(36) := R0 & STA  & '0' & x"11";	-- STA R0, @17	#Constante de limite de valor de minutos e segundos(5)
tmp(37) := R0 & LDI  & '0' & x"03";	-- LDI R0, $3
tmp(38) := R0 & STA  & '0' & x"12";	-- STA R0, @18	#Constante de limite de valor de horas1 (3)
tmp(39) := R0 & LDI  & '0' & x"02";	-- LDI R0, $2
tmp(40) := R0 & STA  & '0' & x"13";	-- STA R0, @19	#Constante de limite de valor de horas2 (2)
tmp(41) := R0 & LDI  & '0' & x"06";	-- LDI R0, $6
tmp(42) := R0 & STA  & '0' & x"14";	-- STA R0, @20	#Constante de limite de valor (6)
tmp(43) := R0 & LDI  & '0' & x"04";	-- LDI R0, $4
tmp(44) := R0 & STA  & '0' & x"15";	-- STA R0, @21	#Constante de limite de valor (4)
tmp(45) := R0 & LDI  & '0' & x"00";	-- LDI R0, $0
tmp(46) := R0 & STA  & '0' & x"16";	-- STA R0, @22	#Flag(0)
tmp(47) := R0 & STA  & '0' & x"1E";	-- STA R0, @30	# Armazena valor para operacao
tmp(48) := R0 & STA  & '0' & x"1F";	-- STA R0, @31
tmp(49) := R0 & STA  & '0' & x"20";	-- STA R0, @32
tmp(50) := R0 & STA  & '0' & x"21";	-- STA R0, @33
tmp(51) := R0 & STA  & '0' & x"22";	-- STA R0, @34
tmp(52) := R0 & STA  & '0' & x"23";	-- STA R0, @35
tmp(53) := R0 & NOP  & '0' & x"00";	-- NOP	#Loop principal
tmp(54) := R2 & LDA  & '1' & x"60";	-- LDA R2, @352	# Le o valor de KEY0
tmp(55) := R2 & CEQ  & '0' & x"06";	-- CEQ R2, @6	# Compara o valor de KEY0 com 0
tmp(56) := R0 & JEQ  & '0' & x"A1";	-- JEQ @PULA1	# Se for igual a 0, nao incrementa e atualiza os displays
tmp(57) := R2 & STA  & '1' & x"FF";	-- STA R2, @511	#Limpa a leitura de KEY0
tmp(58) := R2 & LDA  & '0' & x"00";	-- LDA R2, @0	#Carrega o valor da unidade no acumulador
tmp(59) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na unidade
tmp(60) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara unidade com 10
tmp(61) := R0 & JEQ  & '0' & x"68";	-- JEQ @UNIDADEPASSOU	#Se for igual a 10, incrementa a dezena
tmp(62) := R2 & STA  & '0' & x"00";	-- STA R2, @0	#Se for diferente de 10, armazena o valor da unidade
tmp(63) := R2 & LDA  & '1' & x"61";	-- LDA R2, @353	# Le o valor de KEY1
tmp(64) := R2 & CEQ  & '0' & x"06";	-- CEQ R2, @6	# Compara o valor de KEY1 com 0
tmp(65) := R0 & JEQ  & '0' & x"43";	-- JEQ @CONFEREKEY2	# Se for igual a 0, ignora a subrotina de configuracao de hora
tmp(66) := R0 & JSR  & '0' & x"AF";	-- JSR @CONFIGHORA	# Se for diferente de 0, entra na sub rotina de configuracao de hora
tmp(67) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(68) := R2 & LDA  & '1' & x"62";	-- LDA R2, @354	# Le o valor de KEY2
tmp(69) := R2 & CEQ  & '0' & x"06";	-- CEQ R2, @6	# Compara o valor de KEY2 com 0
tmp(70) := R0 & JEQ  & '0' & x"35";	-- JEQ @INICIOLOOP	# Se for igual a 0, fica no aguardo para quando for 1
tmp(71) := R2 & LDI  & '0' & x"01";	-- LDI R2, $1	# Se for diferente de 0, armazena 1 no acumulador
tmp(72) := R2 & STA  & '0' & x"16";	-- STA R2, @22	#Armazena 1 na flag
tmp(73) := R1 & LDI  & '0' & x"40";	-- LDI R1, $64
tmp(74) := R1 & STA  & '1' & x"00";	-- STA R1, @256
tmp(75) := R2 & LDA  & '0' & x"00";	-- LDA R2, @0
tmp(76) := R2 & STA  & '0' & x"1E";	-- STA R2, @30
tmp(77) := R2 & LDA  & '0' & x"01";	-- LDA R2, @1
tmp(78) := R2 & STA  & '0' & x"1F";	-- STA R2, @31
tmp(79) := R2 & LDA  & '0' & x"02";	-- LDA R2, @2
tmp(80) := R2 & STA  & '0' & x"20";	-- STA R2, @32
tmp(81) := R2 & LDA  & '0' & x"03";	-- LDA R2, @3
tmp(82) := R2 & STA  & '0' & x"21";	-- STA R2, @33
tmp(83) := R2 & LDA  & '0' & x"04";	-- LDA R2, @4
tmp(84) := R2 & STA  & '0' & x"22";	-- STA R2, @34
tmp(85) := R2 & LDA  & '0' & x"05";	-- LDA R2, @5
tmp(86) := R2 & STA  & '0' & x"23";	-- STA R2, @35
tmp(87) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(88) := R2 & LDA  & '0' & x"1E";	-- LDA R2, @30
tmp(89) := R2 & STA  & '0' & x"00";	-- STA R2, @0
tmp(90) := R2 & LDA  & '0' & x"1F";	-- LDA R2, @31
tmp(91) := R2 & STA  & '0' & x"01";	-- STA R2, @1
tmp(92) := R2 & LDA  & '0' & x"20";	-- LDA R2, @32
tmp(93) := R2 & STA  & '0' & x"02";	-- STA R2, @2
tmp(94) := R2 & LDA  & '0' & x"21";	-- LDA R2, @33
tmp(95) := R2 & STA  & '0' & x"03";	-- STA R2, @3
tmp(96) := R2 & LDA  & '0' & x"22";	-- LDA R2, @34
tmp(97) := R2 & STA  & '0' & x"04";	-- STA R2, @4
tmp(98) := R2 & LDA  & '0' & x"23";	-- LDA R2, @35
tmp(99) := R2 & STA  & '0' & x"05";	-- STA R2, @5
tmp(100) := R0 & JSR  & '1' & x"8C";	-- JSR @CHECALIMITE	# Verifica se os valores estao dentro dos limites
tmp(101) := R2 & LDI  & '0' & x"00";	-- LDI R2, $0
tmp(102) := R2 & STA  & '1' & x"00";	-- STA R2, @256
tmp(103) := R0 & JMP  & '0' & x"35";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(104) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(105) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(106) := R2 & STA  & '0' & x"00";	-- STA R2, @0	#Zera a unidade
tmp(107) := R2 & LDA  & '0' & x"01";	-- LDA R2, @1	#Carrega o valor da dezena no acumulador
tmp(108) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na dezena 
tmp(109) := R2 & CEQ  & '0' & x"14";	-- CEQ R2, @20	#Compara dezena com 6
tmp(110) := R2 & JEQ  & '0' & x"71";	-- JEQ R2, @DEZENAPASSOU	#Se for igual a 6, incrementa a centena
tmp(111) := R2 & STA  & '0' & x"01";	-- STA R2, @1	#Se for diferente de 6, armazena o valor da dezena
tmp(112) := R0 & JMP  & '0' & x"35";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(113) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(114) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(115) := R2 & STA  & '0' & x"01";	-- STA R2, @1	#Zera a dezena
tmp(116) := R2 & LDA  & '0' & x"02";	-- LDA R2, @2	#Carrega o valor da centena no acumulador
tmp(117) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na centena
tmp(118) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara centena com 10
tmp(119) := R0 & JEQ  & '0' & x"7A";	-- JEQ @CENTENAPASSOU	#Se for igual a 10, incrementa a unidade de milhar
tmp(120) := R2 & STA  & '0' & x"02";	-- STA R2, @2	#Se for diferente de 10, armazena o valor da centena
tmp(121) := R0 & JMP  & '0' & x"35";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(122) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(123) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(124) := R2 & STA  & '0' & x"02";	-- STA R2, @2	#Zera a centena
tmp(125) := R2 & LDA  & '0' & x"03";	-- LDA R2, @3	#Carrega o valor da unidade de milhar no acumulador
tmp(126) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na unidade de milhar
tmp(127) := R2 & CEQ  & '0' & x"14";	-- CEQ R2, @20	#Compara unidade de milhar com 6
tmp(128) := R0 & JEQ  & '0' & x"83";	-- JEQ @UNIDADEMILHARPASSOU	#Se for igual a 6, incrementa a dezena de milhar
tmp(129) := R2 & STA  & '0' & x"03";	-- STA R2, @3	#Se for diferente de 6, armazena o valor da unidade de milhar
tmp(130) := R0 & JMP  & '0' & x"35";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(131) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(132) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(133) := R2 & STA  & '0' & x"03";	-- STA R2, @3	#Zera a unidade de milhar
tmp(134) := R2 & LDA  & '0' & x"05";	-- LDA R2, @5	#Carrega o valor da centena de milhar no acumulador
tmp(135) := R2 & CEQ  & '0' & x"13";	-- CEQ R2, @19	#Compara com 2
tmp(136) := R0 & JEQ  & '0' & x"8F";	-- JEQ @HORACERTADEZENAMILHAR	#Se for igual a 2, vai pra essa condicao
tmp(137) := R2 & LDA  & '0' & x"04";	-- LDA R2, @4	#Carrega o valor da dezena de milhar no acumulador
tmp(138) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na dezena de milhar
tmp(139) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara dezena de milhar com 10
tmp(140) := R0 & JEQ  & '0' & x"96";	-- JEQ @DEZENAMILHARPASSOU	#Se for igual a 10, incrementa a centena de milhar
tmp(141) := R2 & STA  & '0' & x"04";	-- STA R2, @4	#Se for diferente de 10, armazena o valor da dezena de milhar
tmp(142) := R0 & JMP  & '0' & x"35";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(143) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(144) := R2 & LDA  & '0' & x"04";	-- LDA R2, @4	#Carrega o valor da dezena de milhar no acumulador
tmp(145) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na dezena de milhar
tmp(146) := R2 & CEQ  & '0' & x"15";	-- CEQ R2, @21	#Compara dezena de milhar com 4
tmp(147) := R0 & JEQ  & '0' & x"9F";	-- JEQ @VIROUAHORA	#Se for igual a 4, virou a hora
tmp(148) := R2 & STA  & '0' & x"04";	-- STA R2, @4	#Se for diferente de 4, armazena o valor da dezena de milhar
tmp(149) := R0 & JMP  & '0' & x"35";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(150) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(151) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(152) := R2 & STA  & '0' & x"04";	-- STA R2, @4	#Zera a dezena de milhar
tmp(153) := R2 & LDA  & '0' & x"05";	-- LDA R2, @5	#Carrega o valor da centena de milhar no acumulador
tmp(154) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na centena de milhar
tmp(155) := R2 & CEQ  & '0' & x"12";	-- CEQ R2, @18	#Compara com 3
tmp(156) := R0 & JEQ  & '0' & x"83";	-- JEQ @UNIDADEMILHARPASSOU	#Se for igual a 3, volta
tmp(157) := R2 & STA  & '0' & x"05";	-- STA R2, @5	#Se for diferente de 3, armazena o valor da centena de milhar
tmp(158) := R0 & JMP  & '0' & x"35";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(159) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(160) := R0 & JMP  & '0' & x"00";	-- JMP @RESTART	#Retorna para o LOOP principal
tmp(161) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(162) := R3 & LDA  & '0' & x"00";	-- LDA R3, @0	#Le o valor das unidades
tmp(163) := R3 & STA  & '1' & x"20";	-- STA R3, @288	#Armazena o valor das unidades no HEX0
tmp(164) := R3 & LDA  & '0' & x"01";	-- LDA R3, @1	#Le o valor das dezenas
tmp(165) := R3 & STA  & '1' & x"21";	-- STA R3, @289	#Armazena o valor das dezenas no HEX1
tmp(166) := R3 & LDA  & '0' & x"02";	-- LDA R3, @2	#Le o valor das centenas
tmp(167) := R3 & STA  & '1' & x"22";	-- STA R3, @290	#Armazena o valor das centenas no HEX2
tmp(168) := R3 & LDA  & '0' & x"03";	-- LDA R3, @3	#Le o valor das unidades de milhar
tmp(169) := R3 & STA  & '1' & x"23";	-- STA R3, @291	#Armazena o valor das unidades de milhar no HEX3
tmp(170) := R3 & LDA  & '0' & x"04";	-- LDA R3, @4	#Le o valor das dezenas de milhar
tmp(171) := R3 & STA  & '1' & x"24";	-- STA R3, @292	#Armazena o valor das dezenas de milhar no HEX4
tmp(172) := R3 & LDA  & '0' & x"05";	-- LDA R3, @5	#Le o valor das centenas de milhar
tmp(173) := R3 & STA  & '1' & x"25";	-- STA R3, @293	#Armazena o valor das centenas de milhar no HEX5
tmp(174) := R0 & JMP  & '0' & x"35";	-- JMP @INICIOLOOP	# Volta para o loop principal
tmp(175) := R0 & NOP  & '0' & x"00";	-- NOP	#Rotina de configuracao de hora
tmp(176) := R0 & LDA  & '0' & x"06";	-- LDA R0, @6	#Carrega 0 no acumulador
tmp(177) := R0 & STA  & '0' & x"00";	-- STA R0, @0	#Armazenando 0 em unidade, dezena, centena, etc
tmp(178) := R0 & STA  & '0' & x"01";	-- STA R0, @1
tmp(179) := R0 & STA  & '0' & x"02";	-- STA R0, @2
tmp(180) := R0 & STA  & '0' & x"03";	-- STA R0, @3
tmp(181) := R0 & STA  & '0' & x"04";	-- STA R0, @4
tmp(182) := R0 & STA  & '0' & x"05";	-- STA R0, @5
tmp(183) := R0 & STA  & '1' & x"20";	-- STA R0, @288	# Zera o HEX1
tmp(184) := R0 & STA  & '1' & x"21";	-- STA R0, @289	# Zera o HEX2
tmp(185) := R0 & STA  & '1' & x"22";	-- STA R0, @290	# Zera o HEX3
tmp(186) := R0 & STA  & '1' & x"23";	-- STA R0, @291	# Zera o HEX4
tmp(187) := R0 & STA  & '1' & x"24";	-- STA R0, @292	# Zera o HEX5
tmp(188) := R0 & STA  & '1' & x"25";	-- STA R0, @293	# Zera o HEX6
tmp(189) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1	# Carrega o valor 1
tmp(190) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota no endereco dos LEDS(7-0)
tmp(191) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Limpa a leitura de KEY1
tmp(192) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(193) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(194) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(195) := R0 & JGT  & '0' & x"C5";	-- JGT @VALORATUALIZADO	#Se for maior que 9, atualiza os displays
tmp(196) := R0 & JMP  & '0' & x"C7";	-- JMP @IGNORA
tmp(197) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(198) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(199) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(200) := R1 & STA  & '1' & x"20";	-- STA R1, @288	# Hex 0
tmp(201) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	# Le KEY1
tmp(202) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara KEY1 com 0
tmp(203) := R0 & JEQ  & '0' & x"C0";	-- JEQ @ESPERAUNIDADE	#Se for 0, ou seja, nao esta apertado, espera ate apertar
tmp(204) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Limpa a leitura de KEY1
tmp(205) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(206) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(207) := R0 & JGT  & '0' & x"D1";	-- JGT @VALORATUALIZADO2	#Se for maior que 9, atualiza os displays
tmp(208) := R0 & JMP  & '0' & x"D3";	-- JMP @IGNORA2
tmp(209) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(210) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(211) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(212) := R1 & STA  & '0' & x"00";	-- STA R1, @0	#Armazena o valor das chaves no limite das unidades
tmp(213) := R0 & JMP  & '0' & x"D6";	-- JMP @ESPERADEZENA
tmp(214) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(215) := R1 & LDI  & '0' & x"04";	-- LDI R1, $4	#Carrega o valor 4
tmp(216) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(217) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(218) := R1 & GT  & '0' & x"11";	-- GT R1, @17	#Compara com 5
tmp(219) := R0 & JGT  & '0' & x"DD";	-- JGT @VALORATUALIZADO3	#Se for maior que 5, atualiza os displays
tmp(220) := R0 & JMP  & '0' & x"DF";	-- JMP @IGNORA3
tmp(221) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(222) := R1 & LDI  & '0' & x"05";	-- LDI R1, $5
tmp(223) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(224) := R1 & STA  & '1' & x"21";	-- STA R1, @289	# Hex 1
tmp(225) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(226) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(227) := R0 & JEQ  & '0' & x"D6";	-- JEQ @ESPERADEZENA	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(228) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(229) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(230) := R1 & GT  & '0' & x"11";	-- GT R1, @17	#Compara com 5
tmp(231) := R0 & JGT  & '0' & x"E9";	-- JGT @VALORATUALIZADO4	#Se for maior que 5, atualiza os displays
tmp(232) := R0 & JMP  & '0' & x"EB";	-- JMP @IGNORA4
tmp(233) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(234) := R1 & LDI  & '0' & x"05";	-- LDI R1, $5
tmp(235) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(236) := R1 & STA  & '0' & x"01";	-- STA R1, @1	#Armazena o valor das chaves no limte das dezenas
tmp(237) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(238) := R1 & LDI  & '0' & x"10";	-- LDI R1, $16	# Carrega o valor 16 no acumulador
tmp(239) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(240) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(241) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(242) := R0 & JGT  & '0' & x"F4";	-- JGT @VALORATUALIZADO5	#Se for maior que 9, atualiza os displays
tmp(243) := R0 & JMP  & '0' & x"F6";	-- JMP @IGNORA5
tmp(244) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(245) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(246) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(247) := R1 & STA  & '1' & x"22";	-- STA R1, @290	# Hex 2
tmp(248) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(249) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(250) := R0 & JEQ  & '0' & x"ED";	-- JEQ @ESPERACENTENA	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(251) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(252) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(253) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(254) := R0 & JGT  & '1' & x"00";	-- JGT @VALORATUALIZADO6	#Se for maior que 9, atualiza os displays
tmp(255) := R0 & JMP  & '1' & x"02";	-- JMP @IGNORA6
tmp(256) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(257) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(258) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(259) := R1 & STA  & '0' & x"02";	-- STA R1, @2	#Armazena o valor das chaves no limite das centenas
tmp(260) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(261) := R1 & LDI  & '0' & x"20";	-- LDI R1, $32	# Carrega o valor 32 no acumulador
tmp(262) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(263) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(264) := R1 & GT  & '0' & x"11";	-- GT R1, @17	#Compara com 5
tmp(265) := R0 & JGT  & '1' & x"0B";	-- JGT @VALORATUALIZADO7	#Se for maior que 5, atualiza os displays
tmp(266) := R0 & JMP  & '1' & x"0D";	-- JMP @IGNORA7
tmp(267) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(268) := R1 & LDI  & '0' & x"05";	-- LDI R1, $5
tmp(269) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(270) := R1 & STA  & '1' & x"23";	-- STA R1, @291	# Hex 3
tmp(271) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(272) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1
tmp(273) := R0 & JEQ  & '1' & x"04";	-- JEQ @ESPERAUNIDADEMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(274) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(275) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(276) := R1 & GT  & '0' & x"11";	-- GT R1, @17	#Compara com 5
tmp(277) := R0 & JGT  & '1' & x"17";	-- JGT @VALORATUALIZADO8	#Se for maior que 5, atualiza os displays
tmp(278) := R0 & JMP  & '1' & x"19";	-- JMP @IGNORA8
tmp(279) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(280) := R1 & LDI  & '0' & x"05";	-- LDI R1, $5
tmp(281) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(282) := R1 & STA  & '0' & x"03";	-- STA R1, @3	#Armazena o valor das chaves no limite das unidades de milhar
tmp(283) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(284) := R1 & LDA  & '0' & x"05";	-- LDA R1, @5	#Le o valor da centena de milhar
tmp(285) := R1 & GT  & '0' & x"07";	-- GT R1, @7	#Compara com 1
tmp(286) := R0 & JGT  & '1' & x"36";	-- JGT @AJUSTADEZENAMILHAR
tmp(287) := R1 & LDI  & '0' & x"80";	-- LDI R1, $128	# Carrega o valor 128 no acumulador
tmp(288) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(289) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(290) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(291) := R0 & JGT  & '1' & x"25";	-- JGT @VALORATUALIZADO9	#Se for maior que 9, atualiza os displays
tmp(292) := R0 & JMP  & '1' & x"27";	-- JMP @IGNORA9
tmp(293) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(294) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(295) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(296) := R1 & STA  & '1' & x"24";	-- STA R1, @292	# Hex 4
tmp(297) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(298) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(299) := R0 & JEQ  & '1' & x"1B";	-- JEQ @ESPERADEZENAMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(300) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(301) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(302) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(303) := R0 & JGT  & '1' & x"31";	-- JGT @VALORATUALIZADO10	#Se for maior que 9, atualiza os displays
tmp(304) := R0 & JMP  & '1' & x"33";	-- JMP @IGNORA10
tmp(305) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(306) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(307) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(308) := R1 & STA  & '0' & x"04";	-- STA R1, @4	#Armazena o valor das chaves no limite das dezenas de milhar
tmp(309) := R0 & JMP  & '1' & x"4D";	-- JMP @ESPERACENTENAMILHAR
tmp(310) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(311) := R1 & LDI  & '0' & x"80";	-- LDI R1, $128	# Carrega o valor 128 no acumulador
tmp(312) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(313) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(314) := R1 & GT  & '0' & x"12";	-- GT R1, @18	#Compara com 3
tmp(315) := R0 & JGT  & '1' & x"3D";	-- JGT @VALORATUALIZADO13	#Se for maior que 3, atualiza os displays
tmp(316) := R0 & JMP  & '1' & x"77";	-- JMP @IGNORA13
tmp(317) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(318) := R1 & LDI  & '0' & x"03";	-- LDI R1, $3
tmp(319) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(320) := R1 & STA  & '1' & x"24";	-- STA R1, @292	# Hex 4
tmp(321) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(322) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(323) := R0 & JEQ  & '1' & x"36";	-- JEQ @AJUSTADEZENAMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(324) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(325) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(326) := R1 & GT  & '0' & x"12";	-- GT R1, @18	#Compara com 3
tmp(327) := R0 & JGT  & '1' & x"49";	-- JGT @VALORATUALIZADO14	#Se for maior que 3, atualiza os displays
tmp(328) := R0 & JMP  & '1' & x"83";	-- JMP @IGNORA14
tmp(329) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(330) := R1 & LDI  & '0' & x"03";	-- LDI R1, $3
tmp(331) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(332) := R1 & STA  & '0' & x"04";	-- STA R1, @4	#Armazena o valor das chaves no limite das dezenas de milhar
tmp(333) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(334) := R1 & LDA  & '0' & x"04";	-- LDA R1, @4	#Le o valor da dezena de milhar
tmp(335) := R1 & GT  & '0' & x"12";	-- GT R1, @18	#Compara com 3
tmp(336) := R0 & JGT  & '1' & x"6C";	-- JGT @HORACERTACENTENAMILHAR
tmp(337) := R1 & LDA  & '0' & x"06";	-- LDA R1, @6	#Carrega 0 no acumulador
tmp(338) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Zera o valor nos LEDS(7~0)
tmp(339) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1	# Carrega o valor 1 no acumulador
tmp(340) := R1 & STA  & '1' & x"01";	-- STA R1, @257	# Bota o valor nos LEDS
tmp(341) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(342) := R1 & GT  & '0' & x"13";	-- GT R1, @19	#Compara com 2
tmp(343) := R0 & JGT  & '1' & x"59";	-- JGT @VALORATUALIZADO11	#Se for maior que 2, atualiza os displays
tmp(344) := R0 & JMP  & '1' & x"5B";	-- JMP @IGNORA11
tmp(345) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(346) := R1 & LDI  & '0' & x"02";	-- LDI R1, $2
tmp(347) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(348) := R1 & STA  & '1' & x"25";	-- STA R1, @293	# Hex 5
tmp(349) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(350) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1
tmp(351) := R0 & JEQ  & '1' & x"4D";	-- JEQ @ESPERACENTENAMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(352) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(353) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(354) := R1 & GT  & '0' & x"13";	-- GT R1, @19	#Compara com 2
tmp(355) := R0 & JGT  & '1' & x"65";	-- JGT @VALORATUALIZADO12	#Se for maior que 2, atualiza os displays
tmp(356) := R0 & JMP  & '1' & x"67";	-- JMP @IGNORA12
tmp(357) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(358) := R1 & LDI  & '0' & x"02";	-- LDI R1, $2
tmp(359) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(360) := R1 & STA  & '0' & x"05";	-- STA R1, @5	#Armazena o valor das chaves no limite das centenas de milhar
tmp(361) := R1 & LDI  & '0' & x"00";	-- LDI R1, $0
tmp(362) := R1 & STA  & '1' & x"01";	-- STA R1, @257
tmp(363) := R0 & JMP  & '1' & x"87";	-- JMP @FINALSUB
tmp(364) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(365) := R1 & LDA  & '0' & x"06";	-- LDA R1, @6	#Carrega 0 no acumulador
tmp(366) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Zera o valor nos LEDS(7~0)
tmp(367) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1	# Carrega o valor 1 no acumulador
tmp(368) := R1 & STA  & '1' & x"01";	-- STA R1, @257	# Bota o valor nos LEDS
tmp(369) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(370) := R1 & GT  & '0' & x"07";	-- GT R1, @7	#Compara com 1
tmp(371) := R0 & JGT  & '1' & x"75";	-- JGT @VALORATUALIZADO15	#Se for maior que 1, atualiza os displays
tmp(372) := R0 & JMP  & '1' & x"77";	-- JMP @IGNORA13
tmp(373) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(374) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1
tmp(375) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(376) := R1 & STA  & '1' & x"25";	-- STA R1, @293	# Hex 5
tmp(377) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(378) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1
tmp(379) := R0 & JEQ  & '1' & x"4D";	-- JEQ @ESPERACENTENAMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(380) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(381) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(382) := R1 & GT  & '0' & x"07";	-- GT R1, @7	#Compara com 1
tmp(383) := R0 & JGT  & '1' & x"81";	-- JGT @VALORATUALIZADO16	#Se for maior que 1, atualiza os displays
tmp(384) := R0 & JMP  & '1' & x"83";	-- JMP @IGNORA14
tmp(385) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(386) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1
tmp(387) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(388) := R1 & STA  & '0' & x"05";	-- STA R1, @5	#Armazena o valor das chaves no limite das centenas de milhar
tmp(389) := R1 & LDI  & '0' & x"00";	-- LDI R1, $0
tmp(390) := R1 & STA  & '1' & x"01";	-- STA R1, @257
tmp(391) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(392) := R1 & LDA  & '0' & x"16";	-- LDA R1, @22
tmp(393) := R1 & CEQ  & '0' & x"07";	-- CEQ R1, @7
tmp(394) := R0 & JEQ  & '1' & x"AE";	-- JEQ @TESTE
tmp(395) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(396) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(397) := R1 & LDA  & '0' & x"00";	-- LDA R1, @0	#Le o valor das unidades
tmp(398) := R1 & CEQ  & '0' & x"0A";	-- CEQ R1, @10	#Compara com o valor limite das unidades
tmp(399) := R0 & JEQ  & '1' & x"91";	-- JEQ @CHECADEZENA	#Se for igual, checa se ocorre com as dezenas
tmp(400) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(401) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(402) := R1 & LDA  & '0' & x"01";	-- LDA R1, @1	#Le o valor das dezenas
tmp(403) := R1 & CEQ  & '0' & x"0B";	-- CEQ R1, @11	#Compara com o valor limite das dezenas
tmp(404) := R0 & JEQ  & '1' & x"96";	-- JEQ @CHECACENTENA	#Se for igual, checa se ocorre com as centenas
tmp(405) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(406) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(407) := R1 & LDA  & '0' & x"02";	-- LDA R1, @2	#Le o valor das centenas
tmp(408) := R1 & CEQ  & '0' & x"0C";	-- CEQ R1, @12	#Compara com o valor limite das centenas
tmp(409) := R0 & JEQ  & '1' & x"9B";	-- JEQ @CHECAUNIDADEMILHAR	#Se for igual, checa se ocorre com as unidades de milhar
tmp(410) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(411) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(412) := R1 & LDA  & '0' & x"03";	-- LDA R1, @3	# Le o valor das unidades de milhar
tmp(413) := R1 & CEQ  & '0' & x"0D";	-- CEQ R1, @13	# Compara com o valor limite das unidades de milhar 
tmp(414) := R0 & JEQ  & '1' & x"A0";	-- JEQ @CHECADEZENAMILHAR	#Se for igual, checa se ocorre com as dezenas de milhar
tmp(415) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(416) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(417) := R1 & LDA  & '0' & x"04";	-- LDA R1, @4	# Le o valor das dezenas de milhar
tmp(418) := R1 & CEQ  & '0' & x"0E";	-- CEQ R1, @14	# Compara com o valor limite das dezenas de milhar 
tmp(419) := R0 & JEQ  & '1' & x"A5";	-- JEQ @CHECACENTENAMILHAR	#Se for igual, checa se ocorre com as centenas de milhar
tmp(420) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(421) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(422) := R1 & LDA  & '0' & x"05";	-- LDA R1, @5	# Le o valor das centenas de milhar
tmp(423) := R1 & CEQ  & '0' & x"0F";	-- CEQ R1, @15	# Compara com o valor limite das centenas de milhar 
tmp(424) := R0 & JEQ  & '1' & x"AA";	-- JEQ @BATEUNOLIMITE	#Se for igual, indica que o limite foi batido
tmp(425) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(426) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(427) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1	#Atribui o valor 1 no acumulador
tmp(428) := R1 & STA  & '1' & x"02";	-- STA R1, @258	#Ativa o LED de limite atingido 
tmp(429) := R0 & RET  & '0' & x"00";	-- RET	#Retorna pro LOOP principal
tmp(430) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(431) := R1 & LDA  & '0' & x"00";	-- LDA R1, @0
tmp(432) := R1 & STA  & '0' & x"0A";	-- STA R1, @10
tmp(433) := R1 & LDA  & '0' & x"01";	-- LDA R1, @1
tmp(434) := R1 & STA  & '0' & x"0B";	-- STA R1, @11
tmp(435) := R1 & LDA  & '0' & x"02";	-- LDA R1, @2
tmp(436) := R1 & STA  & '0' & x"0C";	-- STA R1, @12
tmp(437) := R1 & LDA  & '0' & x"03";	-- LDA R1, @3
tmp(438) := R1 & STA  & '0' & x"0D";	-- STA R1, @13
tmp(439) := R1 & LDA  & '0' & x"04";	-- LDA R1, @4
tmp(440) := R1 & STA  & '0' & x"0E";	-- STA R1, @14
tmp(441) := R1 & LDA  & '0' & x"05";	-- LDA R1, @5
tmp(442) := R1 & STA  & '0' & x"0F";	-- STA R1, @15
tmp(443) := R1 & LDI  & '0' & x"00";	-- LDI R1, $0
tmp(444) := R1 & STA  & '0' & x"16";	-- STA R1, @22
tmp(445) := R0 & JMP  & '0' & x"57";	-- JMP @RETORNO





        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;
library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 13;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is
  
  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI	 : std_logic_vector(3 downto 0) := "0100";
  constant STA	 : std_logic_vector(3 downto 0) := "0101";
  constant JMP : std_logic_vector(3 downto 0) := "0110";
  constant JEQ : std_logic_vector(3 downto 0) := "0111";
  constant CEQ : std_logic_vector(3 downto 0) := "1000";
  constant JSR : std_logic_vector(3 downto 0) := "1001";
  constant RET : std_logic_vector(3 downto 0) := "1010";
  constant GT : std_logic_vector(3 downto 0) := "1011";
  constant JGT : std_logic_vector(3 downto 0) := "1100";
  
  constant R0:    std_logic_vector (1 DOWNTO 0)	:= "00";
  constant R1:    std_logic_vector (1 DOWNTO 0)	:= "01";
  constant R2:    std_logic_vector (1 DOWNTO 0)	:= "10";
  constant R3:    std_logic_vector (1 DOWNTO 0)	:= "11";


  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Reset_A, Operacao_ULA
      -- Inicializa os endereços:
tmp(0) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(1) := R0 & LDI  & '0' & x"00";	-- LDI R0, $0	#Início do Setup
tmp(2) := R0 & STA  & '1' & x"20";	-- STA R0, @288	#Zerando hexas
tmp(3) := R0 & STA  & '1' & x"21";	-- STA R0, @289
tmp(4) := R0 & STA  & '1' & x"22";	-- STA R0, @290
tmp(5) := R0 & STA  & '1' & x"23";	-- STA R0, @291
tmp(6) := R0 & STA  & '1' & x"24";	-- STA R0, @292
tmp(7) := R0 & STA  & '1' & x"25";	-- STA R0, @293
tmp(8) := R0 & STA  & '1' & x"00";	-- STA R0, @256	#Zerando leds
tmp(9) := R0 & STA  & '1' & x"01";	-- STA R0, @257
tmp(10) := R0 & STA  & '1' & x"02";	-- STA R0, @258
tmp(11) := R0 & STA  & '0' & x"00";	-- STA R0, @0	#Armazenando 0 em unidade, dezena, centena, etc
tmp(12) := R0 & STA  & '0' & x"01";	-- STA R0, @1
tmp(13) := R0 & STA  & '0' & x"02";	-- STA R0, @2
tmp(14) := R0 & STA  & '0' & x"03";	-- STA R0, @3
tmp(15) := R0 & STA  & '0' & x"04";	-- STA R0, @4
tmp(16) := R0 & STA  & '0' & x"05";	-- STA R0, @5
tmp(17) := R0 & STA  & '0' & x"06";	-- STA R0, @6	#Constante de comparacao (0)
tmp(18) := R0 & STA  & '0' & x"0F";	-- STA R0, @15	#Flag que para contagem
tmp(19) := R0 & STA  & '1' & x"FE";	-- STA R0, @510
tmp(20) := R0 & STA  & '1' & x"FF";	-- STA R0, @511
tmp(21) := R0 & STA  & '1' & x"FD";	-- STA R0, @509
tmp(22) := R0 & LDI  & '0' & x"01";	-- LDI R0, $1
tmp(23) := R0 & STA  & '0' & x"07";	-- STA R0, @7	#Constante de Incremento (1)
tmp(24) := R0 & LDI  & '0' & x"0A";	-- LDI R0, $10
tmp(25) := R0 & STA  & '0' & x"08";	-- STA R0, @8	#Constante de limite no display (10)
tmp(26) := R0 & LDI  & '0' & x"00";	-- LDI R0, $0
tmp(27) := R0 & STA  & '0' & x"09";	-- STA R0, @9	#Limite de contagem em unidade, dezena, centena, etc
tmp(28) := R0 & STA  & '0' & x"0A";	-- STA R0, @10
tmp(29) := R0 & STA  & '0' & x"0B";	-- STA R0, @11
tmp(30) := R0 & STA  & '0' & x"0C";	-- STA R0, @12
tmp(31) := R0 & STA  & '0' & x"0D";	-- STA R0, @13
tmp(32) := R0 & STA  & '0' & x"0E";	-- STA R0, @14
tmp(33) := R0 & LDI  & '0' & x"09";	-- LDI R0, $9
tmp(34) := R0 & STA  & '0' & x"10";	-- STA R0, @16	#Constante de limite de valor
tmp(35) := R0 & LDI  & '0' & x"05";	-- LDI R0, $5
tmp(36) := R0 & STA  & '0' & x"11";	-- STA R0, @17	#Constante de limite de valor de minutos e segundos
tmp(37) := R0 & LDI  & '0' & x"03";	-- LDI R0, $3
tmp(38) := R0 & STA  & '0' & x"12";	-- STA R0, @18	#Constante de limite de valor de horas1 (3)
tmp(39) := R0 & LDI  & '0' & x"02";	-- LDI R0, $2
tmp(40) := R0 & STA  & '0' & x"13";	-- STA R0, @19	#Constante de limite de valor de horas2 (2)
tmp(41) := R0 & LDI  & '0' & x"06";	-- LDI R0, $6
tmp(42) := R0 & STA  & '0' & x"14";	-- STA R0, @20
tmp(43) := R0 & LDI  & '0' & x"04";	-- LDI R0, $4
tmp(44) := R0 & STA  & '0' & x"15";	-- STA R0, @21
tmp(45) := R0 & LDI  & '0' & x"00";	-- LDI R0, $0
tmp(46) := R0 & STA  & '0' & x"16";	-- STA R0, @22
tmp(47) := R0 & NOP  & '0' & x"00";	-- NOP	#Loop principal
tmp(48) := R0 & NOP  & '0' & x"00";	-- NOP	# Incrementa ate chegar no limite de contagem
tmp(49) := R2 & LDA  & '1' & x"60";	-- LDA R2, @352	# Le o valor de KEY0
tmp(50) := R2 & CEQ  & '0' & x"06";	-- CEQ R2, @6	# Compara o valor de KEY0 com 0
tmp(51) := R0 & JEQ  & '0' & x"8A";	-- JEQ @PULA1	# Se for igual a 0, nao incrementa e atualiza os displays
tmp(52) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(53) := R2 & STA  & '1' & x"FF";	-- STA R2, @511	#Limpa a leitura de KEY1
tmp(54) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(55) := R2 & LDA  & '0' & x"00";	-- LDA R2, @0	#Carrega o valor da unidade no acumulador
tmp(56) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na unidade
tmp(57) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara unidade com 10
tmp(58) := R0 & JEQ  & '0' & x"42";	-- JEQ @UNIDADEPASSOU	#Se for igual a 10, incrementa a dezena
tmp(59) := R2 & STA  & '0' & x"00";	-- STA R2, @0	#Se for diferente de 10, armazena o valor da unidade
tmp(60) := R2 & LDA  & '1' & x"61";	-- LDA R2, @353	# Le o valor de KEY1
tmp(61) := R2 & CEQ  & '0' & x"06";	-- CEQ R2, @6	# Compara o valor de KEY1 com 0
tmp(62) := R0 & JEQ  & '0' & x"2F";	-- JEQ @INICIOLOOP	# Se for igual a 0, fica no aguardo para quando for 1
tmp(63) := R0 & JSR  & '0' & x"99";	-- JSR @CONFIGHORA	# Se for diferente de 0, entra na sub rotina de configuracao de hora
tmp(64) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(65) := R0 & JMP  & '0' & x"2F";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(66) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(67) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(68) := R2 & STA  & '0' & x"00";	-- STA R2, @0	#Zera a unidade
tmp(69) := R2 & LDA  & '0' & x"01";	-- LDA R2, @1	#Carrega o valor da dezena no acumulador
tmp(70) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na dezena 
tmp(71) := R2 & CEQ  & '0' & x"14";	-- CEQ R2, @20	#Compara dezena com 6
tmp(72) := R2 & JEQ  & '0' & x"4B";	-- JEQ R2, @DEZENAPASSOU	#Se for igual a 6, incrementa a centena
tmp(73) := R2 & STA  & '0' & x"01";	-- STA R2, @1	#Se for diferente de 6, armazena o valor da dezena
tmp(74) := R0 & JMP  & '0' & x"2F";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(75) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(76) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(77) := R2 & STA  & '0' & x"01";	-- STA R2, @1	#Zera a dezena
tmp(78) := R2 & LDA  & '0' & x"02";	-- LDA R2, @2	#Carrega o valor da centena no acumulador
tmp(79) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na centena
tmp(80) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara centena com 10
tmp(81) := R0 & JEQ  & '0' & x"54";	-- JEQ @CENTENAPASSOU	#Se for igual a 10, incrementa a unidade de milhar
tmp(82) := R2 & STA  & '0' & x"02";	-- STA R2, @2	#Se for diferente de 10, armazena o valor da centena
tmp(83) := R0 & JMP  & '0' & x"2F";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(84) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(85) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(86) := R2 & STA  & '0' & x"02";	-- STA R2, @2	#Zera a centena
tmp(87) := R2 & LDA  & '0' & x"03";	-- LDA R2, @3	#Carrega o valor da unidade de milhar no acumulador
tmp(88) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na unidade de milhar
tmp(89) := R2 & CEQ  & '0' & x"14";	-- CEQ R2, @20	#Compara unidade de milhar com 6
tmp(90) := R0 & JEQ  & '0' & x"5D";	-- JEQ @UNIDADEMILHARPASSOU	#Se for igual a 6, incrementa a dezena de milhar
tmp(91) := R2 & STA  & '0' & x"03";	-- STA R2, @3	#Se for diferente de 6, armazena o valor da unidade de milhar
tmp(92) := R0 & JMP  & '0' & x"2F";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(93) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(94) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(95) := R2 & STA  & '0' & x"03";	-- STA R2, @3	#Zera a unidade de milhar
tmp(96) := R2 & LDA  & '0' & x"05";	-- LDA R2, @5	#Carrega o valor da centena de milhar no acumulador
tmp(97) := R2 & CEQ  & '0' & x"13";	-- CEQ R2, @19	#Compara com 2
tmp(98) := R0 & JEQ  & '0' & x"69";	-- JEQ @HORACERTADEZENAMILHAR	#Se for igual a 2, vai pra essa condicao
tmp(99) := R2 & LDA  & '0' & x"04";	-- LDA R2, @4	#Carrega o valor da dezena de milhar no acumulador
tmp(100) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na dezena de milhar
tmp(101) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara dezena de milhar com 10
tmp(102) := R0 & JEQ  & '0' & x"70";	-- JEQ @DEZENAMILHARPASSOU	#Se for igual a 10, incrementa a centena de milhar
tmp(103) := R2 & STA  & '0' & x"04";	-- STA R2, @4	#Se for diferente de 10, armazena o valor da dezena de milhar
tmp(104) := R0 & JMP  & '0' & x"2F";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(105) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(106) := R2 & LDA  & '0' & x"04";	-- LDA R2, @4	#Carrega o valor da dezena de milhar no acumulador
tmp(107) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na dezena de milhar
tmp(108) := R2 & CEQ  & '0' & x"15";	-- CEQ R2, @21	#Compara dezena de milhar com 4
tmp(109) := R0 & JEQ  & '0' & x"79";	-- JEQ @VIROUAHORA	#Se for igual a 4, virou a hora
tmp(110) := R2 & STA  & '0' & x"04";	-- STA R2, @4	#Se for diferente de 4, armazena o valor da dezena de milhar
tmp(111) := R0 & JMP  & '0' & x"2F";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(112) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(113) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(114) := R2 & STA  & '0' & x"04";	-- STA R2, @4	#Zera a dezena de milhar
tmp(115) := R2 & LDA  & '0' & x"05";	-- LDA R2, @5	#Carrega o valor da centena de milhar no acumulador
tmp(116) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na centena de milhar
tmp(117) := R2 & CEQ  & '0' & x"12";	-- CEQ R2, @18	#Compara com 3
tmp(118) := R0 & JEQ  & '0' & x"5D";	-- JEQ @UNIDADEMILHARPASSOU	#Se for igual a 3, volta
tmp(119) := R2 & STA  & '0' & x"05";	-- STA R2, @5	#Se for diferente de 3, armazena o valor da centena de milhar
tmp(120) := R0 & JMP  & '0' & x"2F";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(121) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(122) := R0 & JSR  & '0' & x"8D";	-- JSR @ZERADISPLAY
tmp(123) := R0 & JMP  & '0' & x"00";	-- JMP @RESTART	#Retorna para o LOOP principal
tmp(124) := R0 & NOP  & '0' & x"00";	-- NOP	#Atualiza os valores dos HEX
tmp(125) := R3 & LDA  & '0' & x"00";	-- LDA R3, @0	#Le o valor das unidades
tmp(126) := R3 & STA  & '1' & x"20";	-- STA R3, @288	#Armazena o valor das unidades no HEX0
tmp(127) := R3 & LDA  & '0' & x"01";	-- LDA R3, @1	#Le o valor das dezenas
tmp(128) := R3 & STA  & '1' & x"21";	-- STA R3, @289	#Armazena o valor das dezenas no HEX1
tmp(129) := R3 & LDA  & '0' & x"02";	-- LDA R3, @2	#Le o valor das centenas
tmp(130) := R3 & STA  & '1' & x"22";	-- STA R3, @290	#Armazena o valor das centenas no HEX2
tmp(131) := R3 & LDA  & '0' & x"03";	-- LDA R3, @3	#Le o valor das unidades de milhar
tmp(132) := R3 & STA  & '1' & x"23";	-- STA R3, @291	#Armazena o valor das unidades de milhar no HEX3
tmp(133) := R3 & LDA  & '0' & x"04";	-- LDA R3, @4	#Le o valor das dezenas de milhar
tmp(134) := R3 & STA  & '1' & x"24";	-- STA R3, @292	#Armazena o valor das dezenas de milhar no HEX4
tmp(135) := R3 & LDA  & '0' & x"05";	-- LDA R3, @5	#Le o valor das centenas de milhar
tmp(136) := R3 & STA  & '1' & x"25";	-- STA R3, @293	#Armazena o valor das centenas de milhar no HEX5
tmp(137) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(138) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(139) := R0 & JSR  & '0' & x"7C";	-- JSR @ATUALIZA	# Atualiza os displays
tmp(140) := R0 & JMP  & '0' & x"30";	-- JMP @INCREMENTADOR	# Volta para o loop principal
tmp(141) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(142) := R0 & LDA  & '0' & x"06";	-- LDA R0, @6	#Carrega 0 no acumulador
tmp(143) := R0 & STA  & '1' & x"20";	-- STA R0, @288	# Zera o HEX1
tmp(144) := R0 & STA  & '1' & x"21";	-- STA R0, @289	# Zera o HEX2
tmp(145) := R0 & STA  & '1' & x"22";	-- STA R0, @290	# Zera o HEX3
tmp(146) := R0 & STA  & '1' & x"23";	-- STA R0, @291	# Zera o HEX4
tmp(147) := R0 & STA  & '1' & x"24";	-- STA R0, @292	# Zera o HEX5
tmp(148) := R0 & STA  & '1' & x"25";	-- STA R0, @293	# Zera o HEX6
tmp(149) := R0 & STA  & '1' & x"00";	-- STA R0, @256	# Zera os LEDS(7~0)
tmp(150) := R0 & STA  & '1' & x"02";	-- STA R0, @258	# Zera os LED(9)
tmp(151) := R0 & STA  & '1' & x"01";	-- STA R0, @257	# Zera os LED(8) 
tmp(152) := R0 & RET  & '0' & x"00";	-- RET
tmp(153) := R0 & NOP  & '0' & x"00";	-- NOP	#Rotina de configuracao de hora
tmp(154) := R0 & LDA  & '0' & x"06";	-- LDA R0, @6	#Carrega 0 no acumulador
tmp(155) := R0 & STA  & '0' & x"00";	-- STA R0, @0	#Armazenando 0 em unidade, dezena, centena, etc
tmp(156) := R0 & STA  & '0' & x"01";	-- STA R0, @1
tmp(157) := R0 & STA  & '0' & x"02";	-- STA R0, @2
tmp(158) := R0 & STA  & '0' & x"03";	-- STA R0, @3
tmp(159) := R0 & STA  & '0' & x"04";	-- STA R0, @4
tmp(160) := R0 & STA  & '0' & x"05";	-- STA R0, @5
tmp(161) := R0 & STA  & '1' & x"20";	-- STA R0, @288	# Zera o HEX1
tmp(162) := R0 & STA  & '1' & x"21";	-- STA R0, @289	# Zera o HEX2
tmp(163) := R0 & STA  & '1' & x"22";	-- STA R0, @290	# Zera o HEX3
tmp(164) := R0 & STA  & '1' & x"23";	-- STA R0, @291	# Zera o HEX4
tmp(165) := R0 & STA  & '1' & x"24";	-- STA R0, @292	# Zera o HEX5
tmp(166) := R0 & STA  & '1' & x"25";	-- STA R0, @293	# Zera o HEX6
tmp(167) := R0 & STA  & '1' & x"00";	-- STA R0, @256	# Zera os LEDS(7~0)
tmp(168) := R0 & STA  & '1' & x"02";	-- STA R0, @258	# Zera os LED(9)
tmp(169) := R0 & STA  & '1' & x"01";	-- STA R0, @257	# Zera os LED(8) 
tmp(170) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1	# Carrega o valor 1
tmp(171) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota no endereco dos LEDS(7-0)
tmp(172) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Limpa a leitura de KEY1
tmp(173) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(174) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(175) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(176) := R0 & JGT  & '0' & x"B2";	-- JGT @VALORATUALIZADO	#Se for maior que 9, atualiza os displays
tmp(177) := R0 & JMP  & '0' & x"B4";	-- JMP @IGNORA
tmp(178) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(179) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(180) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(181) := R1 & STA  & '1' & x"20";	-- STA R1, @288	# Hex 0
tmp(182) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	# Le KEY1
tmp(183) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara KEY1 com 0
tmp(184) := R0 & JEQ  & '0' & x"AD";	-- JEQ @ESPERAUNIDADE	#Se for 0, ou seja, nao esta apertado, espera ate apertar
tmp(185) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Limpa a leitura de KEY1
tmp(186) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(187) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(188) := R0 & JGT  & '0' & x"BE";	-- JGT @VALORATUALIZADO2	#Se for maior que 9, atualiza os displays
tmp(189) := R0 & JMP  & '0' & x"C0";	-- JMP @IGNORA2
tmp(190) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(191) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(192) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(193) := R1 & STA  & '0' & x"00";	-- STA R1, @0	#Armazena o valor das chaves no limite das unidades
tmp(194) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(195) := R1 & LDI  & '0' & x"04";	-- LDI R1, $4	#Carrega o valor 4
tmp(196) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(197) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(198) := R1 & GT  & '0' & x"11";	-- GT R1, @17	#Compara com 5
tmp(199) := R0 & JGT  & '0' & x"C9";	-- JGT @VALORATUALIZADO3	#Se for maior que 5, atualiza os displays
tmp(200) := R0 & JMP  & '0' & x"CB";	-- JMP @IGNORA3
tmp(201) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(202) := R1 & LDI  & '0' & x"05";	-- LDI R1, $5
tmp(203) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(204) := R1 & STA  & '1' & x"21";	-- STA R1, @289	# Hex 1
tmp(205) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(206) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(207) := R0 & JEQ  & '0' & x"C2";	-- JEQ @ESPERADEZENA	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(208) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(209) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(210) := R1 & GT  & '0' & x"11";	-- GT R1, @17	#Compara com 5
tmp(211) := R0 & JGT  & '0' & x"D5";	-- JGT @VALORATUALIZADO4	#Se for maior que 5, atualiza os displays
tmp(212) := R0 & JMP  & '0' & x"D7";	-- JMP @IGNORA4
tmp(213) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(214) := R1 & LDI  & '0' & x"05";	-- LDI R1, $5
tmp(215) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(216) := R1 & STA  & '0' & x"01";	-- STA R1, @1	#Armazena o valor das chaves no limte das dezenas
tmp(217) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(218) := R1 & LDI  & '0' & x"10";	-- LDI R1, $16	# Carrega o valor 16 no acumulador
tmp(219) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(220) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(221) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(222) := R0 & JGT  & '0' & x"E0";	-- JGT @VALORATUALIZADO5	#Se for maior que 9, atualiza os displays
tmp(223) := R0 & JMP  & '0' & x"E2";	-- JMP @IGNORA5
tmp(224) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(225) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(226) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(227) := R1 & STA  & '1' & x"22";	-- STA R1, @290	# Hex 2
tmp(228) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(229) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(230) := R0 & JEQ  & '0' & x"D9";	-- JEQ @ESPERACENTENA	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(231) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(232) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(233) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(234) := R0 & JGT  & '0' & x"EC";	-- JGT @VALORATUALIZADO6	#Se for maior que 9, atualiza os displays
tmp(235) := R0 & JMP  & '0' & x"EE";	-- JMP @IGNORA6
tmp(236) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(237) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(238) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(239) := R1 & STA  & '0' & x"02";	-- STA R1, @2	#Armazena o valor das chaves no limite das centenas
tmp(240) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(241) := R1 & LDI  & '0' & x"20";	-- LDI R1, $32	# Carrega o valor 32 no acumulador
tmp(242) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(243) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(244) := R1 & GT  & '0' & x"11";	-- GT R1, @17	#Compara com 5
tmp(245) := R0 & JGT  & '0' & x"F7";	-- JGT @VALORATUALIZADO7	#Se for maior que 5, atualiza os displays
tmp(246) := R0 & JMP  & '0' & x"F9";	-- JMP @IGNORA7
tmp(247) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(248) := R1 & LDI  & '0' & x"05";	-- LDI R1, $5
tmp(249) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(250) := R1 & STA  & '1' & x"23";	-- STA R1, @291	# Hex 3
tmp(251) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(252) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1
tmp(253) := R0 & JEQ  & '0' & x"F0";	-- JEQ @ESPERAUNIDADEMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(254) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(255) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(256) := R1 & GT  & '0' & x"11";	-- GT R1, @17	#Compara com 5
tmp(257) := R0 & JGT  & '1' & x"03";	-- JGT @VALORATUALIZADO8	#Se for maior que 5, atualiza os displays
tmp(258) := R0 & JMP  & '1' & x"05";	-- JMP @IGNORA8
tmp(259) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(260) := R1 & LDI  & '0' & x"05";	-- LDI R1, $5
tmp(261) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(262) := R1 & STA  & '0' & x"03";	-- STA R1, @3	#Armazena o valor das chaves no limite das unidades de milhar
tmp(263) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(264) := R1 & LDI  & '0' & x"80";	-- LDI R1, $128	# Carrega o valor 128 no acumulador
tmp(265) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(266) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(267) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(268) := R0 & JGT  & '1' & x"0E";	-- JGT @VALORATUALIZADO9	#Se for maior que 9, atualiza os displays
tmp(269) := R0 & JMP  & '1' & x"10";	-- JMP @IGNORA9
tmp(270) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(271) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(272) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(273) := R1 & STA  & '1' & x"24";	-- STA R1, @292	# Hex 4
tmp(274) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(275) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(276) := R0 & JEQ  & '1' & x"07";	-- JEQ @ESPERADEZENAMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(277) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(278) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(279) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(280) := R0 & JGT  & '1' & x"1A";	-- JGT @VALORATUALIZADO10	#Se for maior que 9, atualiza os displays
tmp(281) := R0 & JMP  & '1' & x"1C";	-- JMP @IGNORA10
tmp(282) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(283) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(284) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(285) := R1 & STA  & '0' & x"04";	-- STA R1, @4	#Armazena o valor das chaves no limite das dezenas de milhar
tmp(286) := R0 & JMP  & '1' & x"36";	-- JMP @ESPERACENTENAMILHAR
tmp(287) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(288) := R1 & LDI  & '0' & x"80";	-- LDI R1, $128	# Carrega o valor 128 no acumulador
tmp(289) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(290) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(291) := R1 & GT  & '0' & x"12";	-- GT R1, @18	#Compara com 3
tmp(292) := R0 & JGT  & '1' & x"26";	-- JGT @VALORATUALIZADO13	#Se for maior que 3, atualiza os displays
tmp(293) := R0 & JMP  & '1' & x"28";	-- JMP @IGNORA13
tmp(294) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(295) := R1 & LDI  & '0' & x"03";	-- LDI R1, $3
tmp(296) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(297) := R1 & STA  & '1' & x"24";	-- STA R1, @292	# Hex 4
tmp(298) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(299) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(300) := R0 & JEQ  & '1' & x"1F";	-- JEQ @VOLTADEZENAMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(301) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(302) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(303) := R1 & GT  & '0' & x"12";	-- GT R1, @18	#Compara com 3
tmp(304) := R0 & JGT  & '1' & x"32";	-- JGT @VALORATUALIZADO14	#Se for maior que 3, atualiza os displays
tmp(305) := R0 & JMP  & '1' & x"34";	-- JMP @IGNORA14
tmp(306) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(307) := R1 & LDI  & '0' & x"03";	-- LDI R1, $3
tmp(308) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(309) := R1 & STA  & '0' & x"04";	-- STA R1, @4	#Armazena o valor das chaves no limite das dezenas de milhar
tmp(310) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(311) := R1 & LDA  & '0' & x"06";	-- LDA R1, @6	#Carrega 0 no acumulador
tmp(312) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Zera o valor nos LEDS(7~0)
tmp(313) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1	# Carrega o valor 1 no acumulador
tmp(314) := R1 & STA  & '1' & x"01";	-- STA R1, @257	# Bota o valor nos LEDS
tmp(315) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(316) := R1 & GT  & '0' & x"13";	-- GT R1, @19	#Compara com 2
tmp(317) := R0 & JGT  & '1' & x"3F";	-- JGT @VALORATUALIZADO11	#Se for maior que 2, atualiza os displays
tmp(318) := R0 & JMP  & '1' & x"41";	-- JMP @IGNORA11
tmp(319) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(320) := R1 & LDI  & '0' & x"02";	-- LDI R1, $2
tmp(321) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(322) := R1 & STA  & '1' & x"25";	-- STA R1, @293	# Hex 5
tmp(323) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(324) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1
tmp(325) := R0 & JEQ  & '1' & x"36";	-- JEQ @ESPERACENTENAMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(326) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(327) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(328) := R1 & GT  & '0' & x"13";	-- GT R1, @19	#Compara com 2
tmp(329) := R0 & JGT  & '1' & x"4B";	-- JGT @VALORATUALIZADO12	#Se for maior que 2, atualiza os displays
tmp(330) := R0 & JMP  & '1' & x"4D";	-- JMP @IGNORA12
tmp(331) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(332) := R1 & LDI  & '0' & x"02";	-- LDI R1, $2
tmp(333) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(334) := R1 & STA  & '0' & x"05";	-- STA R1, @5	#Armazena o valor das chaves no limite das centenas de milhar
tmp(335) := R1 & LDA  & '0' & x"05";	-- LDA R1, @5
tmp(336) := R1 & SOMA  & '0' & x"04";	-- SOMA R1, @4
tmp(337) := R1 & GT  & '0' & x"14";	-- GT R1, @20
tmp(338) := R0 & JGT  & '1' & x"1F";	-- JGT @VOLTADEZENAMILHAR
tmp(339) := R1 & LDI  & '0' & x"00";	-- LDI R1, $0
tmp(340) := R1 & STA  & '1' & x"01";	-- STA R1, @257
tmp(341) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal

        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;
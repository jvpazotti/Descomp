library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 13;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is
  
  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI	 : std_logic_vector(3 downto 0) := "0100";
  constant STA	 : std_logic_vector(3 downto 0) := "0101";
  constant JMP : std_logic_vector(3 downto 0) := "0110";
  constant JEQ : std_logic_vector(3 downto 0) := "0111";
  constant CEQ : std_logic_vector(3 downto 0) := "1000";
  constant JSR : std_logic_vector(3 downto 0) := "1001";
  constant RET : std_logic_vector(3 downto 0) := "1010";
  constant GT : std_logic_vector(3 downto 0) := "1011";
  constant JGT : std_logic_vector(3 downto 0) := "1100";
  
  constant R0:    std_logic_vector (1 DOWNTO 0)	:= "00";
  constant R1:    std_logic_vector (1 DOWNTO 0)	:= "01";
  constant R2:    std_logic_vector (1 DOWNTO 0)	:= "10";
  constant R3:    std_logic_vector (1 DOWNTO 0)	:= "11";


  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Reset_A, Operacao_ULA
      -- Inicializa os endereços:
tmp(0) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(1) := R0 & LDI  & '0' & x"00";	-- LDI R0, $0	#Início do Setup
tmp(2) := R0 & STA  & '1' & x"20";	-- STA R0, @288	#Zerando hexas
tmp(3) := R0 & STA  & '1' & x"21";	-- STA R0, @289
tmp(4) := R0 & STA  & '1' & x"22";	-- STA R0, @290
tmp(5) := R0 & STA  & '1' & x"23";	-- STA R0, @291
tmp(6) := R0 & STA  & '1' & x"24";	-- STA R0, @292
tmp(7) := R0 & STA  & '1' & x"25";	-- STA R0, @293
tmp(8) := R0 & STA  & '1' & x"00";	-- STA R0, @256	#Zerando leds
tmp(9) := R0 & STA  & '1' & x"01";	-- STA R0, @257
tmp(10) := R0 & STA  & '1' & x"02";	-- STA R0, @258
tmp(11) := R0 & STA  & '0' & x"00";	-- STA R0, @0	#Armazenando 0 em unidade, dezena, centena, etc
tmp(12) := R0 & STA  & '0' & x"01";	-- STA R0, @1
tmp(13) := R0 & STA  & '0' & x"02";	-- STA R0, @2
tmp(14) := R0 & STA  & '0' & x"03";	-- STA R0, @3
tmp(15) := R0 & STA  & '0' & x"04";	-- STA R0, @4
tmp(16) := R0 & STA  & '0' & x"05";	-- STA R0, @5
tmp(17) := R0 & STA  & '0' & x"06";	-- STA R0, @6	#Constante de comparacao (0)
tmp(18) := R0 & STA  & '0' & x"0F";	-- STA R0, @15	#Flag que para contagem
tmp(19) := R0 & STA  & '1' & x"FE";	-- STA R0, @510
tmp(20) := R0 & STA  & '1' & x"FF";	-- STA R0, @511
tmp(21) := R0 & STA  & '1' & x"FD";	-- STA R0, @509
tmp(22) := R0 & LDI  & '0' & x"01";	-- LDI R0, $1
tmp(23) := R0 & STA  & '0' & x"07";	-- STA R0, @7	#Constante de Incremento (1)
tmp(24) := R0 & LDI  & '0' & x"0A";	-- LDI R0, $10
tmp(25) := R0 & STA  & '0' & x"08";	-- STA R0, @8	#Constante de limite no display (10)
tmp(26) := R0 & LDI  & '0' & x"00";	-- LDI R0, $0
tmp(27) := R0 & STA  & '0' & x"09";	-- STA R0, @9	#Limite de contagem em unidade, dezena, centena, etc
tmp(28) := R0 & STA  & '0' & x"0A";	-- STA R0, @10
tmp(29) := R0 & STA  & '0' & x"0B";	-- STA R0, @11
tmp(30) := R0 & STA  & '0' & x"0C";	-- STA R0, @12
tmp(31) := R0 & STA  & '0' & x"0D";	-- STA R0, @13
tmp(32) := R0 & STA  & '0' & x"0E";	-- STA R0, @14
tmp(33) := R0 & LDI  & '0' & x"09";	-- LDI R0, $9
tmp(34) := R0 & STA  & '0' & x"10";	-- STA R0, @16	#Constante de limite de valor
tmp(35) := R0 & NOP  & '0' & x"00";	-- NOP	#Loop principal
tmp(36) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	# Le o valor de KEY1
tmp(37) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	# Compara o valor de KEY1 com 0
tmp(38) := R0 & JEQ  & '0' & x"23";	-- JEQ @INICIOLOOP	# Se for igual a 0, fica no aguardo para quando for 1
tmp(39) := R0 & JSR  & '0' & x"3E";	-- JSR @CONFIGLIMITE	# Se for diferente de 0, entra na sub rotina de configuracao de Limite
tmp(40) := R0 & LDA  & '0' & x"06";	-- LDA R0, @6	#Carrega 0 no acumulador
tmp(41) := R0 & STA  & '1' & x"20";	-- STA R0, @288	# Zera o HEX1
tmp(42) := R0 & STA  & '1' & x"21";	-- STA R0, @289	# Zera o HEX2
tmp(43) := R0 & STA  & '1' & x"22";	-- STA R0, @290	# Zera o HEX3
tmp(44) := R0 & STA  & '1' & x"23";	-- STA R0, @291	# Zera o HEX4
tmp(45) := R0 & STA  & '1' & x"24";	-- STA R0, @292	# Zera o HEX5
tmp(46) := R0 & STA  & '1' & x"25";	-- STA R0, @293	# Zera o HEX6
tmp(47) := R0 & STA  & '1' & x"00";	-- STA R0, @256	# Zera os LEDS(7~0)
tmp(48) := R0 & STA  & '1' & x"02";	-- STA R0, @258	# Zera os LED(9)
tmp(49) := R0 & STA  & '1' & x"01";	-- STA R0, @257	# Zera os LED(8) 
tmp(50) := R0 & NOP  & '0' & x"00";	-- NOP	# Incrementa ate chegar no limite de contagem
tmp(51) := R2 & LDA  & '1' & x"60";	-- LDA R2, @352	# Le o valor de KEY0
tmp(52) := R2 & CEQ  & '0' & x"06";	-- CEQ R2, @6	# Compara o valor de KEY0 com 0
tmp(53) := R0 & JEQ  & '0' & x"37";	-- JEQ @PULA1	# Se for igual a 0, nao incrementa e atualiza os displays
tmp(54) := R0 & JSR  & '0' & x"CD";	-- JSR @INCREMENTA	# Se for diferente de 0, entra na sub rotina de incremento
tmp(55) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(56) := R0 & JSR  & '1' & x"0A";	-- JSR @ATUALIZA	# Atualiza os displays
tmp(57) := R0 & JSR  & '1' & x"18";	-- JSR @CHECALIMITE	# Checa pra ver se passou do limite setado
tmp(58) := R2 & LDA  & '0' & x"0F";	-- LDA R2, @15	# Le o valor da flag de inibir contagem
tmp(59) := R2 & CEQ  & '0' & x"06";	-- CEQ R2, @6	# Compara com 0 a flag (flag com valor 1 -> ativa, flag com valor 0 -> desativada)
tmp(60) := R0 & JEQ  & '0' & x"32";	-- JEQ @INCREMENTADOR	#Se a flag for 0, pode continuar incrementando
tmp(61) := R0 & JMP  & '1' & x"3B";	-- JMP @TRAVA	# Se for 1, trava a contagem
tmp(62) := R0 & NOP  & '0' & x"00";	-- NOP	#Rotina de configuracao de limite
tmp(63) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1	# Carrega o valor 1
tmp(64) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota no endereco dos LEDS(7-0)
tmp(65) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Limpa a leitura de KEY1
tmp(66) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(67) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(68) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(69) := R0 & JGT  & '0' & x"47";	-- JGT @VALORATUALIZADO	#Se for maior que 9, atualiza os displays
tmp(70) := R0 & JMP  & '0' & x"49";	-- JMP @IGNORA
tmp(71) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(72) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(73) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(74) := R1 & STA  & '1' & x"20";	-- STA R1, @288	# Hex 0
tmp(75) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	# Le KEY1
tmp(76) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara KEY1 com 0
tmp(77) := R0 & JEQ  & '0' & x"42";	-- JEQ @ESPERAUNIDADE	#Se for 0, ou seja, nao esta apertado, espera ate apertar
tmp(78) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Limpa a leitura de KEY1
tmp(79) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(80) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(81) := R0 & JGT  & '0' & x"53";	-- JGT @VALORATUALIZADO2	#Se for maior que 9, atualiza os displays
tmp(82) := R0 & JMP  & '0' & x"55";	-- JMP @IGNORA2
tmp(83) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(84) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(85) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(86) := R1 & STA  & '0' & x"09";	-- STA R1, @9	#Armazena o valor das chaves no limite das unidades
tmp(87) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(88) := R1 & LDI  & '0' & x"04";	-- LDI R1, $4	#Carrega o valor 4
tmp(89) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(90) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(91) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(92) := R0 & JGT  & '0' & x"5E";	-- JGT @VALORATUALIZADO3	#Se for maior que 9, atualiza os displays
tmp(93) := R0 & JMP  & '0' & x"60";	-- JMP @IGNORA3
tmp(94) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(95) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(96) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(97) := R1 & STA  & '1' & x"21";	-- STA R1, @289	# Hex 1
tmp(98) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(99) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(100) := R0 & JEQ  & '0' & x"57";	-- JEQ @ESPERADEZENA	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(101) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(102) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(103) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(104) := R0 & JGT  & '0' & x"6A";	-- JGT @VALORATUALIZADO4	#Se for maior que 9, atualiza os displays
tmp(105) := R0 & JMP  & '0' & x"6C";	-- JMP @IGNORA4
tmp(106) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(107) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(108) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(109) := R1 & STA  & '0' & x"0A";	-- STA R1, @10	#Armazena o valor das chaves no limte das dezenas
tmp(110) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(111) := R1 & LDI  & '0' & x"10";	-- LDI R1, $16	# Carrega o valor 16 no acumulador
tmp(112) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(113) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(114) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(115) := R0 & JGT  & '0' & x"75";	-- JGT @VALORATUALIZADO5	#Se for maior que 9, atualiza os displays
tmp(116) := R0 & JMP  & '0' & x"77";	-- JMP @IGNORA5
tmp(117) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(118) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(119) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(120) := R1 & STA  & '1' & x"22";	-- STA R1, @290	# Hex 2
tmp(121) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(122) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(123) := R0 & JEQ  & '0' & x"6E";	-- JEQ @ESPERACENTENA	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(124) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(125) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(126) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(127) := R0 & JGT  & '0' & x"81";	-- JGT @VALORATUALIZADO6	#Se for maior que 9, atualiza os displays
tmp(128) := R0 & JMP  & '0' & x"83";	-- JMP @IGNORA6
tmp(129) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(130) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(131) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(132) := R1 & STA  & '0' & x"0B";	-- STA R1, @11	#Armazena o valor das chaves no limite das centenas
tmp(133) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(134) := R1 & LDI  & '0' & x"20";	-- LDI R1, $32	# Carrega o valor 32 no acumulador
tmp(135) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(136) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(137) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(138) := R0 & JGT  & '0' & x"8C";	-- JGT @VALORATUALIZADO7	#Se for maior que 9, atualiza os displays
tmp(139) := R0 & JMP  & '0' & x"8E";	-- JMP @IGNORA7
tmp(140) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(141) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(142) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(143) := R1 & STA  & '1' & x"23";	-- STA R1, @291	# Hex 3
tmp(144) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(145) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1
tmp(146) := R0 & JEQ  & '0' & x"85";	-- JEQ @ESPERAUNIDADEMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(147) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(148) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(149) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(150) := R0 & JGT  & '0' & x"98";	-- JGT @VALORATUALIZADO8	#Se for maior que 9, atualiza os displays
tmp(151) := R0 & JMP  & '0' & x"9A";	-- JMP @IGNORA8
tmp(152) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(153) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(154) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(155) := R1 & STA  & '0' & x"0C";	-- STA R1, @12	#Armazena o valor das chaves no limite das unidades de milhar
tmp(156) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(157) := R1 & LDI  & '0' & x"80";	-- LDI R1, $128	# Carrega o valor 128 no acumulador
tmp(158) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(159) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(160) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(161) := R0 & JGT  & '0' & x"A3";	-- JGT @VALORATUALIZADO9	#Se for maior que 9, atualiza os displays
tmp(162) := R0 & JMP  & '0' & x"A5";	-- JMP @IGNORA9
tmp(163) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(164) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(165) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(166) := R1 & STA  & '1' & x"24";	-- STA R1, @292	# Hex 4
tmp(167) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(168) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(169) := R0 & JEQ  & '0' & x"9C";	-- JEQ @ESPERADEZENAMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(170) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(171) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(172) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(173) := R0 & JGT  & '0' & x"AF";	-- JGT @VALORATUALIZADO10	#Se for maior que 9, atualiza os displays
tmp(174) := R0 & JMP  & '0' & x"B1";	-- JMP @IGNORA10
tmp(175) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(176) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(177) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(178) := R1 & STA  & '0' & x"0D";	-- STA R1, @13	#Armazena o valor das chaves no limite das dezenas de milhar
tmp(179) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(180) := R1 & LDA  & '0' & x"06";	-- LDA R1, @6	#Carrega 0 no acumulador
tmp(181) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Zera o valor nos LEDS(7~0)
tmp(182) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1	# Carrega o valor 1 no acumulador
tmp(183) := R1 & STA  & '1' & x"01";	-- STA R1, @257	# Bota o valor nos LEDS
tmp(184) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(185) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(186) := R0 & JGT  & '0' & x"BC";	-- JGT @VALORATUALIZADO11	#Se for maior que 9, atualiza os displays
tmp(187) := R0 & JMP  & '0' & x"BE";	-- JMP @IGNORA11
tmp(188) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(189) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(190) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(191) := R1 & STA  & '1' & x"25";	-- STA R1, @293	# Hex 5
tmp(192) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(193) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1
tmp(194) := R0 & JEQ  & '0' & x"B3";	-- JEQ @ESPERACENTENAMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(195) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(196) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(197) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(198) := R0 & JGT  & '0' & x"C8";	-- JGT @VALORATUALIZADO12	#Se for maior que 9, atualiza os displays
tmp(199) := R0 & JMP  & '0' & x"CA";	-- JMP @IGNORA12
tmp(200) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(201) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(202) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(203) := R1 & STA  & '0' & x"0E";	-- STA R1, @14	#Armazena o valor das chaves no limite das centenas de milhar
tmp(204) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(205) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(206) := R2 & STA  & '1' & x"FF";	-- STA R2, @511	#Limpa a leitura de KEY1
tmp(207) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(208) := R2 & LDA  & '0' & x"00";	-- LDA R2, @0	#Carrega o valor da unidade no acumulador
tmp(209) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na unidade
tmp(210) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara unidade com 10
tmp(211) := R0 & JEQ  & '0' & x"D6";	-- JEQ @UNIDADEPASSOU	#Se for igual a 10, incrementa a dezena
tmp(212) := R2 & STA  & '0' & x"00";	-- STA R2, @0	#Se for diferente de 10, armazena o valor da unidade
tmp(213) := R0 & RET  & '0' & x"00";	-- RET 	#Retorna para o LOOP principal
tmp(214) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(215) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(216) := R2 & STA  & '0' & x"00";	-- STA R2, @0	#Zera a unidade
tmp(217) := R2 & LDA  & '0' & x"01";	-- LDA R2, @1	#Carrega o valor da dezena no acumulador
tmp(218) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na dezena 
tmp(219) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara dezena com 10
tmp(220) := R2 & JEQ  & '0' & x"DF";	-- JEQ R2, @DEZENAPASSOU	#Se for igual a 10, incrementa a centena
tmp(221) := R2 & STA  & '0' & x"01";	-- STA R2, @1	#Se for diferente de 10, armazena o valor da dezena
tmp(222) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(223) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(224) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(225) := R2 & STA  & '0' & x"01";	-- STA R2, @1	#Zera a dezena
tmp(226) := R2 & LDA  & '0' & x"02";	-- LDA R2, @2	#Carrega o valor da centena no acumulador
tmp(227) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na centena
tmp(228) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara centena com 10
tmp(229) := R0 & JEQ  & '0' & x"E8";	-- JEQ @CENTENAPASSOU	#Se for igual a 10, incrementa a unidade de milhar
tmp(230) := R2 & STA  & '0' & x"02";	-- STA R2, @2	#Se for diferente de 10, armazena o valor da centena
tmp(231) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(232) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(233) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(234) := R2 & STA  & '0' & x"02";	-- STA R2, @2	#Zera a centena
tmp(235) := R2 & LDA  & '0' & x"03";	-- LDA R2, @3	#Carrega o valor da unidade de milhar no acumulador
tmp(236) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na unidade de milhar
tmp(237) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara unidade de milhar com 10
tmp(238) := R0 & JEQ  & '0' & x"F1";	-- JEQ @UNIDADEMILHARPASSOU	#Se for igual a 10, incrementa a dezena de milhar
tmp(239) := R2 & STA  & '0' & x"03";	-- STA R2, @3	#Se for diferente de 10, armazena o valor da unidade de milhar
tmp(240) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(241) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(242) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(243) := R2 & STA  & '0' & x"03";	-- STA R2, @3	#Zera a unidade de milhar
tmp(244) := R2 & LDA  & '0' & x"04";	-- LDA R2, @4	#Carrega o valor da dezena de milhar no acumulador
tmp(245) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na dezena de milhar
tmp(246) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara dezena de milhar com 10
tmp(247) := R0 & JEQ  & '0' & x"FA";	-- JEQ @DEZENAMILHARPASSOU	#Se for igual a 10, incrementa a centena de milhar
tmp(248) := R2 & STA  & '0' & x"04";	-- STA R2, @4	#Se for diferente de 10, armazena o valor da dezena de milhar
tmp(249) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(250) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(251) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(252) := R2 & STA  & '0' & x"04";	-- STA R2, @4	#Zera a dezena de milhar
tmp(253) := R2 & LDA  & '0' & x"05";	-- LDA R2, @5	#Carrega o valor da centena de milhar no acumulador
tmp(254) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na centena de milhar
tmp(255) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara centena de milhar com 10
tmp(256) := R0 & JEQ  & '1' & x"03";	-- JEQ @CENTENAMILHARPASSOU	#Se for igual a 10, incrementa a unidade de milhao
tmp(257) := R2 & STA  & '0' & x"05";	-- STA R2, @5	#Se for diferente de 10, armazena o valor da centena de milhar
tmp(258) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(259) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(260) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(261) := R2 & STA  & '0' & x"05";	-- STA R2, @5	#Zera a centena de milhar
tmp(262) := R2 & LDI  & '0' & x"01";	-- LDI R2, $1	#Carrega 1 no acumulador
tmp(263) := R2 & STA  & '1' & x"02";	-- STA R2, @258	#Acende o LED(9)
tmp(264) := R2 & STA  & '0' & x"0F";	-- STA R2, @15	#Ativa a flag de inibir incremento
tmp(265) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(266) := R0 & NOP  & '0' & x"00";	-- NOP	#Atualiza os valores dos HEX
tmp(267) := R3 & LDA  & '0' & x"00";	-- LDA R3, @0	#Le o valor das unidades
tmp(268) := R3 & STA  & '1' & x"20";	-- STA R3, @288	#Armazena o valor das unidades no HEX0
tmp(269) := R3 & LDA  & '0' & x"01";	-- LDA R3, @1	#Le o valor das dezenas
tmp(270) := R3 & STA  & '1' & x"21";	-- STA R3, @289	#Armazena o valor das dezenas no HEX1
tmp(271) := R3 & LDA  & '0' & x"02";	-- LDA R3, @2	#Le o valor das centenas
tmp(272) := R3 & STA  & '1' & x"22";	-- STA R3, @290	#Armazena o valor das centenas no HEX2
tmp(273) := R3 & LDA  & '0' & x"03";	-- LDA R3, @3	#Le o valor das unidades de milhar
tmp(274) := R3 & STA  & '1' & x"23";	-- STA R3, @291	#Armazena o valor das unidades de milhar no HEX3
tmp(275) := R3 & LDA  & '0' & x"04";	-- LDA R3, @4	#Le o valor das dezenas de milhar
tmp(276) := R3 & STA  & '1' & x"24";	-- STA R3, @292	#Armazena o valor das dezenas de milhar no HEX4
tmp(277) := R3 & LDA  & '0' & x"05";	-- LDA R3, @5	#Le o valor das centenas de milhar
tmp(278) := R3 & STA  & '1' & x"25";	-- STA R3, @293	#Armazena o valor das centenas de milhar no HEX5
tmp(279) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(280) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(281) := R1 & LDA  & '0' & x"00";	-- LDA R1, @0	#Le o valor das unidades
tmp(282) := R1 & CEQ  & '0' & x"09";	-- CEQ R1, @9	#Compara com o valor limite das unidades
tmp(283) := R0 & JEQ  & '1' & x"1D";	-- JEQ @CHECADEZENA	#Se for igual, checa se ocorre com as dezenas
tmp(284) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(285) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(286) := R1 & LDA  & '0' & x"01";	-- LDA R1, @1	#Le o valor das dezenas
tmp(287) := R1 & CEQ  & '0' & x"0A";	-- CEQ R1, @10	#Compara com o valor limite das dezenas
tmp(288) := R0 & JEQ  & '1' & x"22";	-- JEQ @CHECACENTENA	#Se for igual, checa se ocorre com as centenas
tmp(289) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(290) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(291) := R1 & LDA  & '0' & x"02";	-- LDA R1, @2	#Le o valor das centenas
tmp(292) := R1 & CEQ  & '0' & x"0B";	-- CEQ R1, @11	#Compara com o valor limite das centenas
tmp(293) := R0 & JEQ  & '1' & x"27";	-- JEQ @CHECAUNIDADEMILHAR	#Se for igual, checa se ocorre com as unidades de milhar
tmp(294) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(295) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(296) := R1 & LDA  & '0' & x"03";	-- LDA R1, @3	# Le o valor das unidades de milhar
tmp(297) := R1 & CEQ  & '0' & x"0C";	-- CEQ R1, @12	# Compara com o valor limite das unidades de milhar 
tmp(298) := R0 & JEQ  & '1' & x"2C";	-- JEQ @CHECADEZENAMILHAR	#Se for igual, checa se ocorre com as dezenas de milhar
tmp(299) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(300) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(301) := R1 & LDA  & '0' & x"04";	-- LDA R1, @4	# Le o valor das dezenas de milhar
tmp(302) := R1 & CEQ  & '0' & x"0D";	-- CEQ R1, @13	# Compara com o valor limite das dezenas de milhar 
tmp(303) := R0 & JEQ  & '1' & x"31";	-- JEQ @CHECACENTENAMILHAR	#Se for igual, checa se ocorre com as centenas de milhar
tmp(304) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(305) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(306) := R1 & LDA  & '0' & x"05";	-- LDA R1, @5	# Le o valor das centenas de milhar
tmp(307) := R1 & CEQ  & '0' & x"0E";	-- CEQ R1, @14	# Compara com o valor limite das centenas de milhar 
tmp(308) := R0 & JEQ  & '1' & x"36";	-- JEQ @BATEUNOLIMITE	#Se for igual, indica que o limite foi batido
tmp(309) := R0 & RET  & '0' & x"00";	-- RET	#Se for diferente, retorna para o LOOP principal
tmp(310) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(311) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1	#Atribui o valor 1 no acumulador
tmp(312) := R1 & STA  & '0' & x"0F";	-- STA R1, @15	#Ativa a flag de parar contagem
tmp(313) := R1 & STA  & '1' & x"02";	-- STA R1, @258	#Ativa o LED de limite atingido 
tmp(314) := R0 & RET  & '0' & x"00";	-- RET	#Retorna pro LOOP principal
tmp(315) := R0 & NOP  & '0' & x"00";	-- NOP	#Trava a contagem
tmp(316) := R3 & LDI  & '0' & x"01";	-- LDI R3, $1
tmp(317) := R3 & STA  & '1' & x"00";	-- STA R3, @256
tmp(318) := R3 & LDA  & '1' & x"64";	-- LDA R3, @356	#Le o valor do botao FPGA
tmp(319) := R3 & CEQ  & '0' & x"06";	-- CEQ R3, @6	#Compara com 0 o botao FPGA
tmp(320) := R0 & JEQ  & '1' & x"3B";	-- JEQ @TRAVA	#Se for igual, continua travado
tmp(321) := R0 & JMP  & '0' & x"00";	-- JMP @RESTART	#Se for diferente, reinicia a contagem





        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;
library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 13;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is
  
  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI	 : std_logic_vector(3 downto 0) := "0100";
  constant STA	 : std_logic_vector(3 downto 0) := "0101";
  constant JMP : std_logic_vector(3 downto 0) := "0110";
  constant JEQ : std_logic_vector(3 downto 0) := "0111";
  constant CEQ : std_logic_vector(3 downto 0) := "1000";
  constant JSR : std_logic_vector(3 downto 0) := "1001";
  constant RET : std_logic_vector(3 downto 0) := "1010";
  constant GT : std_logic_vector(3 downto 0) := "1011";
  constant JGT : std_logic_vector(3 downto 0) := "1100";
  
  constant R0:    std_logic_vector (1 DOWNTO 0)	:= "00";
  constant R1:    std_logic_vector (1 DOWNTO 0)	:= "01";
  constant R2:    std_logic_vector (1 DOWNTO 0)	:= "10";
  constant R3:    std_logic_vector (1 DOWNTO 0)	:= "11";


  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Reset_A, Operacao_ULA
      -- Inicializa os endereços:
tmp(0) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(1) := R0 & LDI  & '0' & x"00";	-- LDI R0, $0	#Início do Setup
tmp(2) := R0 & STA  & '1' & x"20";	-- STA R0, @288	#Zerando hexas
tmp(3) := R0 & STA  & '1' & x"21";	-- STA R0, @289
tmp(4) := R0 & STA  & '1' & x"22";	-- STA R0, @290
tmp(5) := R0 & STA  & '1' & x"23";	-- STA R0, @291
tmp(6) := R0 & STA  & '1' & x"24";	-- STA R0, @292
tmp(7) := R0 & STA  & '1' & x"25";	-- STA R0, @293
tmp(8) := R0 & STA  & '1' & x"00";	-- STA R0, @256	#Zerando leds
tmp(9) := R0 & STA  & '1' & x"01";	-- STA R0, @257
tmp(10) := R0 & STA  & '1' & x"02";	-- STA R0, @258
tmp(11) := R0 & STA  & '0' & x"00";	-- STA R0, @0	#Armazenando 0 em unidade, dezena, centena, etc
tmp(12) := R0 & STA  & '0' & x"01";	-- STA R0, @1
tmp(13) := R0 & STA  & '0' & x"02";	-- STA R0, @2
tmp(14) := R0 & STA  & '0' & x"03";	-- STA R0, @3
tmp(15) := R0 & STA  & '0' & x"04";	-- STA R0, @4
tmp(16) := R0 & STA  & '0' & x"05";	-- STA R0, @5
tmp(17) := R0 & STA  & '0' & x"06";	-- STA R0, @6	#Constante de comparacao (0)
tmp(18) := R0 & STA  & '1' & x"FE";	-- STA R0, @510
tmp(19) := R0 & STA  & '1' & x"FF";	-- STA R0, @511
tmp(20) := R0 & STA  & '1' & x"FD";	-- STA R0, @509
tmp(21) := R0 & LDI  & '0' & x"01";	-- LDI R0, $1
tmp(22) := R0 & STA  & '0' & x"07";	-- STA R0, @7	#Constante de Incremento (1)
tmp(23) := R0 & LDI  & '0' & x"0A";	-- LDI R0, $10
tmp(24) := R0 & STA  & '0' & x"08";	-- STA R0, @8	#Constante de limite no display (10)
tmp(25) := R0 & LDI  & '0' & x"00";	-- LDI R0, $0
tmp(26) := R0 & STA  & '0' & x"09";	-- STA R0, @9	#Limite de contagem em unidade, dezena, centena, etc
tmp(27) := R0 & STA  & '0' & x"0A";	-- STA R0, @10
tmp(28) := R0 & STA  & '0' & x"0B";	-- STA R0, @11
tmp(29) := R0 & STA  & '0' & x"0C";	-- STA R0, @12
tmp(30) := R0 & STA  & '0' & x"0D";	-- STA R0, @13
tmp(31) := R0 & STA  & '0' & x"0E";	-- STA R0, @14
tmp(32) := R0 & STA  & '0' & x"0F";	-- STA R0, @15
tmp(33) := R0 & LDI  & '0' & x"09";	-- LDI R0, $9
tmp(34) := R0 & STA  & '0' & x"10";	-- STA R0, @16	#Constante de limite de valor(9)
tmp(35) := R0 & LDI  & '0' & x"05";	-- LDI R0, $5
tmp(36) := R0 & STA  & '0' & x"11";	-- STA R0, @17	#Constante de limite de valor de minutos e segundos(5)
tmp(37) := R0 & LDI  & '0' & x"03";	-- LDI R0, $3
tmp(38) := R0 & STA  & '0' & x"12";	-- STA R0, @18	#Constante de limite de valor de horas1 (3)
tmp(39) := R0 & LDI  & '0' & x"02";	-- LDI R0, $2
tmp(40) := R0 & STA  & '0' & x"13";	-- STA R0, @19	#Constante de limite de valor de horas2 (2)
tmp(41) := R0 & LDI  & '0' & x"06";	-- LDI R0, $6
tmp(42) := R0 & STA  & '0' & x"14";	-- STA R0, @20	#Constante de limite de valor (6)
tmp(43) := R0 & LDI  & '0' & x"04";	-- LDI R0, $4
tmp(44) := R0 & STA  & '0' & x"15";	-- STA R0, @21	#Constante de limite de valor (4)
tmp(45) := R0 & LDI  & '0' & x"00";	-- LDI R0, $0
tmp(46) := R0 & STA  & '0' & x"16";	-- STA R0, @22	#Flag(0)
tmp(47) := R0 & NOP  & '0' & x"00";	-- NOP	#Loop principal
tmp(48) := R2 & LDA  & '1' & x"60";	-- LDA R2, @352	# Le o valor de KEY0
tmp(49) := R2 & CEQ  & '0' & x"06";	-- CEQ R2, @6	# Compara o valor de KEY0 com 0
tmp(50) := R0 & JEQ  & '0' & x"8C";	-- JEQ @PULA1	# Se for igual a 0, nao incrementa e atualiza os displays
tmp(51) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(52) := R2 & STA  & '1' & x"FF";	-- STA R2, @511	#Limpa a leitura de KEY1
tmp(53) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(54) := R2 & LDA  & '0' & x"00";	-- LDA R2, @0	#Carrega o valor da unidade no acumulador
tmp(55) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na unidade
tmp(56) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara unidade com 10
tmp(57) := R0 & JEQ  & '0' & x"45";	-- JEQ @UNIDADEPASSOU	#Se for igual a 10, incrementa a dezena
tmp(58) := R2 & STA  & '0' & x"00";	-- STA R2, @0	#Se for diferente de 10, armazena o valor da unidade
tmp(59) := R2 & LDA  & '1' & x"61";	-- LDA R2, @353	# Le o valor de KEY1
tmp(60) := R2 & CEQ  & '0' & x"06";	-- CEQ R2, @6	# Compara o valor de KEY1 com 0
tmp(61) := R0 & JEQ  & '0' & x"3F";	-- JEQ @CONFEREKEY2	# Se for igual a 0, ignora a subrotina de configuracao de hora
tmp(62) := R0 & JSR  & '0' & x"8F";	-- JSR @CONFIGHORA	# Se for diferente de 0, entra na sub rotina de configuracao de hora
tmp(63) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(64) := R2 & LDA  & '1' & x"62";	-- LDA R2, @354	# Le o valor de KEY2
tmp(65) := R2 & CEQ  & '0' & x"06";	-- CEQ R2, @6	# Compara o valor de KEY2 com 0
tmp(66) := R0 & JEQ  & '0' & x"2F";	-- JEQ @INICIOLOOP	# Se for igual a 0, fica no aguardo para quando for 1
tmp(67) := R0 & JSR  & '1' & x"6B";	-- JSR @ALARME	# Se for diferente de 0, entra na sub rotina de configuracao de alarme
tmp(68) := R0 & JMP  & '0' & x"2F";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(69) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(70) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(71) := R2 & STA  & '0' & x"00";	-- STA R2, @0	#Zera a unidade
tmp(72) := R2 & LDA  & '0' & x"01";	-- LDA R2, @1	#Carrega o valor da dezena no acumulador
tmp(73) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na dezena 
tmp(74) := R2 & CEQ  & '0' & x"14";	-- CEQ R2, @20	#Compara dezena com 6
tmp(75) := R2 & JEQ  & '0' & x"4E";	-- JEQ R2, @DEZENAPASSOU	#Se for igual a 6, incrementa a centena
tmp(76) := R2 & STA  & '0' & x"01";	-- STA R2, @1	#Se for diferente de 6, armazena o valor da dezena
tmp(77) := R0 & JMP  & '0' & x"2F";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(78) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(79) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(80) := R2 & STA  & '0' & x"01";	-- STA R2, @1	#Zera a dezena
tmp(81) := R2 & LDA  & '0' & x"02";	-- LDA R2, @2	#Carrega o valor da centena no acumulador
tmp(82) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na centena
tmp(83) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara centena com 10
tmp(84) := R0 & JEQ  & '0' & x"57";	-- JEQ @CENTENAPASSOU	#Se for igual a 10, incrementa a unidade de milhar
tmp(85) := R2 & STA  & '0' & x"02";	-- STA R2, @2	#Se for diferente de 10, armazena o valor da centena
tmp(86) := R0 & JMP  & '0' & x"2F";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(87) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(88) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(89) := R2 & STA  & '0' & x"02";	-- STA R2, @2	#Zera a centena
tmp(90) := R2 & LDA  & '0' & x"03";	-- LDA R2, @3	#Carrega o valor da unidade de milhar no acumulador
tmp(91) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na unidade de milhar
tmp(92) := R2 & CEQ  & '0' & x"14";	-- CEQ R2, @20	#Compara unidade de milhar com 6
tmp(93) := R0 & JEQ  & '0' & x"60";	-- JEQ @UNIDADEMILHARPASSOU	#Se for igual a 6, incrementa a dezena de milhar
tmp(94) := R2 & STA  & '0' & x"03";	-- STA R2, @3	#Se for diferente de 6, armazena o valor da unidade de milhar
tmp(95) := R0 & JMP  & '0' & x"2F";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(96) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(97) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(98) := R2 & STA  & '0' & x"03";	-- STA R2, @3	#Zera a unidade de milhar
tmp(99) := R2 & LDA  & '0' & x"05";	-- LDA R2, @5	#Carrega o valor da centena de milhar no acumulador
tmp(100) := R2 & CEQ  & '0' & x"13";	-- CEQ R2, @19	#Compara com 2
tmp(101) := R0 & JEQ  & '0' & x"6C";	-- JEQ @HORACERTADEZENAMILHAR	#Se for igual a 2, vai pra essa condicao
tmp(102) := R2 & LDA  & '0' & x"04";	-- LDA R2, @4	#Carrega o valor da dezena de milhar no acumulador
tmp(103) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na dezena de milhar
tmp(104) := R2 & CEQ  & '0' & x"08";	-- CEQ R2, @8	#Compara dezena de milhar com 10
tmp(105) := R0 & JEQ  & '0' & x"73";	-- JEQ @DEZENAMILHARPASSOU	#Se for igual a 10, incrementa a centena de milhar
tmp(106) := R2 & STA  & '0' & x"04";	-- STA R2, @4	#Se for diferente de 10, armazena o valor da dezena de milhar
tmp(107) := R0 & JMP  & '0' & x"2F";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(108) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(109) := R2 & LDA  & '0' & x"04";	-- LDA R2, @4	#Carrega o valor da dezena de milhar no acumulador
tmp(110) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na dezena de milhar
tmp(111) := R2 & CEQ  & '0' & x"15";	-- CEQ R2, @21	#Compara dezena de milhar com 4
tmp(112) := R0 & JEQ  & '0' & x"7C";	-- JEQ @VIROUAHORA	#Se for igual a 4, virou a hora
tmp(113) := R2 & STA  & '0' & x"04";	-- STA R2, @4	#Se for diferente de 4, armazena o valor da dezena de milhar
tmp(114) := R0 & JMP  & '0' & x"2F";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(115) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(116) := R2 & LDA  & '0' & x"06";	-- LDA R2, @6	#Carrega 0 no acumulador
tmp(117) := R2 & STA  & '0' & x"04";	-- STA R2, @4	#Zera a dezena de milhar
tmp(118) := R2 & LDA  & '0' & x"05";	-- LDA R2, @5	#Carrega o valor da centena de milhar no acumulador
tmp(119) := R2 & SOMA  & '0' & x"07";	-- SOMA R2, @7	#Incrementa 1 na centena de milhar
tmp(120) := R2 & CEQ  & '0' & x"12";	-- CEQ R2, @18	#Compara com 3
tmp(121) := R0 & JEQ  & '0' & x"60";	-- JEQ @UNIDADEMILHARPASSOU	#Se for igual a 3, volta
tmp(122) := R2 & STA  & '0' & x"05";	-- STA R2, @5	#Se for diferente de 3, armazena o valor da centena de milhar
tmp(123) := R0 & JMP  & '0' & x"2F";	-- JMP @INICIOLOOP	#Retorna para o LOOP principal
tmp(124) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(125) := R0 & JMP  & '0' & x"00";	-- JMP @RESTART	#Retorna para o LOOP principal
tmp(126) := R0 & NOP  & '0' & x"00";	-- NOP	#Atualiza os valores dos HEX
tmp(127) := R3 & LDA  & '0' & x"00";	-- LDA R3, @0	#Le o valor das unidades
tmp(128) := R3 & STA  & '1' & x"20";	-- STA R3, @288	#Armazena o valor das unidades no HEX0
tmp(129) := R3 & LDA  & '0' & x"01";	-- LDA R3, @1	#Le o valor das dezenas
tmp(130) := R3 & STA  & '1' & x"21";	-- STA R3, @289	#Armazena o valor das dezenas no HEX1
tmp(131) := R3 & LDA  & '0' & x"02";	-- LDA R3, @2	#Le o valor das centenas
tmp(132) := R3 & STA  & '1' & x"22";	-- STA R3, @290	#Armazena o valor das centenas no HEX2
tmp(133) := R3 & LDA  & '0' & x"03";	-- LDA R3, @3	#Le o valor das unidades de milhar
tmp(134) := R3 & STA  & '1' & x"23";	-- STA R3, @291	#Armazena o valor das unidades de milhar no HEX3
tmp(135) := R3 & LDA  & '0' & x"04";	-- LDA R3, @4	#Le o valor das dezenas de milhar
tmp(136) := R3 & STA  & '1' & x"24";	-- STA R3, @292	#Armazena o valor das dezenas de milhar no HEX4
tmp(137) := R3 & LDA  & '0' & x"05";	-- LDA R3, @5	#Le o valor das centenas de milhar
tmp(138) := R3 & STA  & '1' & x"25";	-- STA R3, @293	#Armazena o valor das centenas de milhar no HEX5
tmp(139) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(140) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(141) := R0 & JSR  & '0' & x"7E";	-- JSR @ATUALIZA	# Atualiza os displays
tmp(142) := R0 & JMP  & '0' & x"2F";	-- JMP @INICIOLOOP	# Volta para o loop principal
tmp(143) := R0 & NOP  & '0' & x"00";	-- NOP	#Rotina de configuracao de hora
tmp(144) := R0 & LDA  & '0' & x"06";	-- LDA R0, @6	#Carrega 0 no acumulador
tmp(145) := R0 & STA  & '0' & x"00";	-- STA R0, @0	#Armazenando 0 em unidade, dezena, centena, etc
tmp(146) := R0 & STA  & '0' & x"01";	-- STA R0, @1
tmp(147) := R0 & STA  & '0' & x"02";	-- STA R0, @2
tmp(148) := R0 & STA  & '0' & x"03";	-- STA R0, @3
tmp(149) := R0 & STA  & '0' & x"04";	-- STA R0, @4
tmp(150) := R0 & STA  & '0' & x"05";	-- STA R0, @5
tmp(151) := R0 & STA  & '1' & x"20";	-- STA R0, @288	# Zera o HEX1
tmp(152) := R0 & STA  & '1' & x"21";	-- STA R0, @289	# Zera o HEX2
tmp(153) := R0 & STA  & '1' & x"22";	-- STA R0, @290	# Zera o HEX3
tmp(154) := R0 & STA  & '1' & x"23";	-- STA R0, @291	# Zera o HEX4
tmp(155) := R0 & STA  & '1' & x"24";	-- STA R0, @292	# Zera o HEX5
tmp(156) := R0 & STA  & '1' & x"25";	-- STA R0, @293	# Zera o HEX6
tmp(157) := R0 & STA  & '1' & x"00";	-- STA R0, @256	# Zera os LEDS(7~0)
tmp(158) := R0 & STA  & '1' & x"02";	-- STA R0, @258	# Zera os LED(9)
tmp(159) := R0 & STA  & '1' & x"01";	-- STA R0, @257	# Zera os LED(8) 
tmp(160) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1	# Carrega o valor 1
tmp(161) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota no endereco dos LEDS(7-0)
tmp(162) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Limpa a leitura de KEY1
tmp(163) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(164) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(165) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(166) := R0 & JGT  & '0' & x"A8";	-- JGT @VALORATUALIZADO	#Se for maior que 9, atualiza os displays
tmp(167) := R0 & JMP  & '0' & x"AA";	-- JMP @IGNORA
tmp(168) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(169) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(170) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(171) := R1 & STA  & '1' & x"20";	-- STA R1, @288	# Hex 0
tmp(172) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	# Le KEY1
tmp(173) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara KEY1 com 0
tmp(174) := R0 & JEQ  & '0' & x"A3";	-- JEQ @ESPERAUNIDADE	#Se for 0, ou seja, nao esta apertado, espera ate apertar
tmp(175) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Limpa a leitura de KEY1
tmp(176) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(177) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(178) := R0 & JGT  & '0' & x"B4";	-- JGT @VALORATUALIZADO2	#Se for maior que 9, atualiza os displays
tmp(179) := R0 & JMP  & '0' & x"B6";	-- JMP @IGNORA2
tmp(180) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(181) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(182) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(183) := R1 & STA  & '0' & x"00";	-- STA R1, @0	#Armazena o valor das chaves no limite das unidades
tmp(184) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(185) := R1 & LDI  & '0' & x"04";	-- LDI R1, $4	#Carrega o valor 4
tmp(186) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(187) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(188) := R1 & GT  & '0' & x"11";	-- GT R1, @17	#Compara com 5
tmp(189) := R0 & JGT  & '0' & x"BF";	-- JGT @VALORATUALIZADO3	#Se for maior que 5, atualiza os displays
tmp(190) := R0 & JMP  & '0' & x"C1";	-- JMP @IGNORA3
tmp(191) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(192) := R1 & LDI  & '0' & x"05";	-- LDI R1, $5
tmp(193) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(194) := R1 & STA  & '1' & x"21";	-- STA R1, @289	# Hex 1
tmp(195) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(196) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(197) := R0 & JEQ  & '0' & x"B8";	-- JEQ @ESPERADEZENA	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(198) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(199) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(200) := R1 & GT  & '0' & x"11";	-- GT R1, @17	#Compara com 5
tmp(201) := R0 & JGT  & '0' & x"CB";	-- JGT @VALORATUALIZADO4	#Se for maior que 5, atualiza os displays
tmp(202) := R0 & JMP  & '0' & x"CD";	-- JMP @IGNORA4
tmp(203) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(204) := R1 & LDI  & '0' & x"05";	-- LDI R1, $5
tmp(205) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(206) := R1 & STA  & '0' & x"01";	-- STA R1, @1	#Armazena o valor das chaves no limte das dezenas
tmp(207) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(208) := R1 & LDI  & '0' & x"10";	-- LDI R1, $16	# Carrega o valor 16 no acumulador
tmp(209) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(210) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(211) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(212) := R0 & JGT  & '0' & x"D6";	-- JGT @VALORATUALIZADO5	#Se for maior que 9, atualiza os displays
tmp(213) := R0 & JMP  & '0' & x"D8";	-- JMP @IGNORA5
tmp(214) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(215) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(216) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(217) := R1 & STA  & '1' & x"22";	-- STA R1, @290	# Hex 2
tmp(218) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(219) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(220) := R0 & JEQ  & '0' & x"CF";	-- JEQ @ESPERACENTENA	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(221) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(222) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(223) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(224) := R0 & JGT  & '0' & x"E2";	-- JGT @VALORATUALIZADO6	#Se for maior que 9, atualiza os displays
tmp(225) := R0 & JMP  & '0' & x"E4";	-- JMP @IGNORA6
tmp(226) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(227) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(228) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(229) := R1 & STA  & '0' & x"02";	-- STA R1, @2	#Armazena o valor das chaves no limite das centenas
tmp(230) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(231) := R1 & LDI  & '0' & x"20";	-- LDI R1, $32	# Carrega o valor 32 no acumulador
tmp(232) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(233) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(234) := R1 & GT  & '0' & x"11";	-- GT R1, @17	#Compara com 5
tmp(235) := R0 & JGT  & '0' & x"ED";	-- JGT @VALORATUALIZADO7	#Se for maior que 5, atualiza os displays
tmp(236) := R0 & JMP  & '0' & x"EF";	-- JMP @IGNORA7
tmp(237) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(238) := R1 & LDI  & '0' & x"05";	-- LDI R1, $5
tmp(239) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(240) := R1 & STA  & '1' & x"23";	-- STA R1, @291	# Hex 3
tmp(241) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(242) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1
tmp(243) := R0 & JEQ  & '0' & x"E6";	-- JEQ @ESPERAUNIDADEMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(244) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(245) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(246) := R1 & GT  & '0' & x"11";	-- GT R1, @17	#Compara com 5
tmp(247) := R0 & JGT  & '0' & x"F9";	-- JGT @VALORATUALIZADO8	#Se for maior que 5, atualiza os displays
tmp(248) := R0 & JMP  & '0' & x"FB";	-- JMP @IGNORA8
tmp(249) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(250) := R1 & LDI  & '0' & x"05";	-- LDI R1, $5
tmp(251) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(252) := R1 & STA  & '0' & x"03";	-- STA R1, @3	#Armazena o valor das chaves no limite das unidades de milhar
tmp(253) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(254) := R1 & LDA  & '0' & x"05";	-- LDA R1, @5	#Le o valor da centena de milhar
tmp(255) := R1 & GT  & '0' & x"07";	-- GT R1, @7	#Compara com 1
tmp(256) := R0 & JGT  & '1' & x"18";	-- JGT @AJUSTADEZENAMILHAR
tmp(257) := R1 & LDI  & '0' & x"80";	-- LDI R1, $128	# Carrega o valor 128 no acumulador
tmp(258) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(259) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(260) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(261) := R0 & JGT  & '1' & x"07";	-- JGT @VALORATUALIZADO9	#Se for maior que 9, atualiza os displays
tmp(262) := R0 & JMP  & '1' & x"09";	-- JMP @IGNORA9
tmp(263) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(264) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(265) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(266) := R1 & STA  & '1' & x"24";	-- STA R1, @292	# Hex 4
tmp(267) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(268) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(269) := R0 & JEQ  & '0' & x"FD";	-- JEQ @ESPERADEZENAMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(270) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(271) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(272) := R1 & GT  & '0' & x"10";	-- GT R1, @16	#Compara com 9
tmp(273) := R0 & JGT  & '1' & x"13";	-- JGT @VALORATUALIZADO10	#Se for maior que 9, atualiza os displays
tmp(274) := R0 & JMP  & '1' & x"15";	-- JMP @IGNORA10
tmp(275) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(276) := R1 & LDI  & '0' & x"09";	-- LDI R1, $9
tmp(277) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(278) := R1 & STA  & '0' & x"04";	-- STA R1, @4	#Armazena o valor das chaves no limite das dezenas de milhar
tmp(279) := R0 & JMP  & '1' & x"2F";	-- JMP @ESPERACENTENAMILHAR
tmp(280) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(281) := R1 & LDI  & '0' & x"80";	-- LDI R1, $128	# Carrega o valor 128 no acumulador
tmp(282) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Bota o valor nos LEDS
tmp(283) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(284) := R1 & GT  & '0' & x"12";	-- GT R1, @18	#Compara com 3
tmp(285) := R0 & JGT  & '1' & x"1F";	-- JGT @VALORATUALIZADO13	#Se for maior que 3, atualiza os displays
tmp(286) := R0 & JMP  & '1' & x"59";	-- JMP @IGNORA13
tmp(287) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(288) := R1 & LDI  & '0' & x"03";	-- LDI R1, $3
tmp(289) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(290) := R1 & STA  & '1' & x"24";	-- STA R1, @292	# Hex 4
tmp(291) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(292) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1 
tmp(293) := R0 & JEQ  & '1' & x"18";	-- JEQ @AJUSTADEZENAMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(294) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(295) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(296) := R1 & GT  & '0' & x"12";	-- GT R1, @18	#Compara com 3
tmp(297) := R0 & JGT  & '1' & x"2B";	-- JGT @VALORATUALIZADO14	#Se for maior que 3, atualiza os displays
tmp(298) := R0 & JMP  & '1' & x"65";	-- JMP @IGNORA14
tmp(299) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(300) := R1 & LDI  & '0' & x"03";	-- LDI R1, $3
tmp(301) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(302) := R1 & STA  & '0' & x"04";	-- STA R1, @4	#Armazena o valor das chaves no limite das dezenas de milhar
tmp(303) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(304) := R1 & LDA  & '0' & x"04";	-- LDA R1, @4	#Le o valor da dezena de milhar
tmp(305) := R1 & GT  & '0' & x"12";	-- GT R1, @18	#Compara com 3
tmp(306) := R0 & JGT  & '1' & x"4E";	-- JGT @HORACERTACENTENAMILHAR
tmp(307) := R1 & LDA  & '0' & x"06";	-- LDA R1, @6	#Carrega 0 no acumulador
tmp(308) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Zera o valor nos LEDS(7~0)
tmp(309) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1	# Carrega o valor 1 no acumulador
tmp(310) := R1 & STA  & '1' & x"01";	-- STA R1, @257	# Bota o valor nos LEDS
tmp(311) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(312) := R1 & GT  & '0' & x"13";	-- GT R1, @19	#Compara com 2
tmp(313) := R0 & JGT  & '1' & x"3B";	-- JGT @VALORATUALIZADO11	#Se for maior que 2, atualiza os displays
tmp(314) := R0 & JMP  & '1' & x"3D";	-- JMP @IGNORA11
tmp(315) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(316) := R1 & LDI  & '0' & x"02";	-- LDI R1, $2
tmp(317) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(318) := R1 & STA  & '1' & x"25";	-- STA R1, @293	# Hex 5
tmp(319) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(320) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1
tmp(321) := R0 & JEQ  & '1' & x"2F";	-- JEQ @ESPERACENTENAMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(322) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(323) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(324) := R1 & GT  & '0' & x"13";	-- GT R1, @19	#Compara com 2
tmp(325) := R0 & JGT  & '1' & x"47";	-- JGT @VALORATUALIZADO12	#Se for maior que 2, atualiza os displays
tmp(326) := R0 & JMP  & '1' & x"49";	-- JMP @IGNORA12
tmp(327) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(328) := R1 & LDI  & '0' & x"02";	-- LDI R1, $2
tmp(329) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(330) := R1 & STA  & '0' & x"05";	-- STA R1, @5	#Armazena o valor das chaves no limite das centenas de milhar
tmp(331) := R1 & LDI  & '0' & x"00";	-- LDI R1, $0
tmp(332) := R1 & STA  & '1' & x"01";	-- STA R1, @257
tmp(333) := R0 & JMP  & '1' & x"69";	-- JMP @FINALSUB
tmp(334) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(335) := R1 & LDA  & '0' & x"06";	-- LDA R1, @6	#Carrega 0 no acumulador
tmp(336) := R1 & STA  & '1' & x"00";	-- STA R1, @256	# Zera o valor nos LEDS(7~0)
tmp(337) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1	# Carrega o valor 1 no acumulador
tmp(338) := R1 & STA  & '1' & x"01";	-- STA R1, @257	# Bota o valor nos LEDS
tmp(339) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(340) := R1 & GT  & '0' & x"07";	-- GT R1, @7	#Compara com 1
tmp(341) := R0 & JGT  & '1' & x"57";	-- JGT @VALORATUALIZADO15	#Se for maior que 1, atualiza os displays
tmp(342) := R0 & JMP  & '1' & x"59";	-- JMP @IGNORA13
tmp(343) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(344) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1
tmp(345) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(346) := R1 & STA  & '1' & x"25";	-- STA R1, @293	# Hex 5
tmp(347) := R1 & LDA  & '1' & x"61";	-- LDA R1, @353	#Le o valor de KEY1 novamente
tmp(348) := R1 & CEQ  & '0' & x"06";	-- CEQ R1, @6	#Compara com 0 o valor de KEY1
tmp(349) := R0 & JEQ  & '1' & x"2F";	-- JEQ @ESPERACENTENAMILHAR	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(350) := R1 & STA  & '1' & x"FE";	-- STA R1, @510	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(351) := R1 & LDA  & '1' & x"40";	-- LDA R1, @320	#Le o valor das chaves SW(7~0)
tmp(352) := R1 & GT  & '0' & x"07";	-- GT R1, @7	#Compara com 1
tmp(353) := R0 & JGT  & '1' & x"63";	-- JGT @VALORATUALIZADO16	#Se for maior que 1, atualiza os displays
tmp(354) := R0 & JMP  & '1' & x"65";	-- JMP @IGNORA14
tmp(355) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(356) := R1 & LDI  & '0' & x"01";	-- LDI R1, $1
tmp(357) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(358) := R1 & STA  & '0' & x"05";	-- STA R1, @5	#Armazena o valor das chaves no limite das centenas de milhar
tmp(359) := R1 & LDI  & '0' & x"00";	-- LDI R1, $0
tmp(360) := R1 & STA  & '1' & x"01";	-- STA R1, @257
tmp(361) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(362) := R0 & RET  & '0' & x"00";	-- RET	#Retorna para o LOOP principal
tmp(363) := R0 & NOP  & '0' & x"00";	-- NOP
tmp(364) := R0 & RET  & '0' & x"00";	-- RET



        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;